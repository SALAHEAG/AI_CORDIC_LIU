magic
tech sky130A
magscale 1 2
timestamp 1695408310
<< obsli1 >>
rect 1104 2159 18860 47345
<< obsm1 >>
rect 14 2128 19766 47376
<< metal2 >>
rect 202 49200 258 50000
rect 570 49200 626 50000
rect 1030 49200 1086 50000
rect 1398 49200 1454 50000
rect 1858 49200 1914 50000
rect 2318 49200 2374 50000
rect 2686 49200 2742 50000
rect 3146 49200 3202 50000
rect 3514 49200 3570 50000
rect 3974 49200 4030 50000
rect 4434 49200 4490 50000
rect 4802 49200 4858 50000
rect 5262 49200 5318 50000
rect 5722 49200 5778 50000
rect 6090 49200 6146 50000
rect 6550 49200 6606 50000
rect 6918 49200 6974 50000
rect 7378 49200 7434 50000
rect 7838 49200 7894 50000
rect 8206 49200 8262 50000
rect 8666 49200 8722 50000
rect 9034 49200 9090 50000
rect 9494 49200 9550 50000
rect 9954 49200 10010 50000
rect 10322 49200 10378 50000
rect 10782 49200 10838 50000
rect 11242 49200 11298 50000
rect 11610 49200 11666 50000
rect 12070 49200 12126 50000
rect 12438 49200 12494 50000
rect 12898 49200 12954 50000
rect 13358 49200 13414 50000
rect 13726 49200 13782 50000
rect 14186 49200 14242 50000
rect 14554 49200 14610 50000
rect 15014 49200 15070 50000
rect 15474 49200 15530 50000
rect 15842 49200 15898 50000
rect 16302 49200 16358 50000
rect 16762 49200 16818 50000
rect 17130 49200 17186 50000
rect 17590 49200 17646 50000
rect 17958 49200 18014 50000
rect 18418 49200 18474 50000
rect 18878 49200 18934 50000
rect 19246 49200 19302 50000
rect 19706 49200 19762 50000
rect 1398 0 1454 800
rect 4250 0 4306 800
rect 7102 0 7158 800
rect 9954 0 10010 800
rect 12806 0 12862 800
rect 15658 0 15714 800
rect 18510 0 18566 800
<< obsm2 >>
rect 20 49144 146 49314
rect 314 49144 514 49314
rect 682 49144 974 49314
rect 1142 49144 1342 49314
rect 1510 49144 1802 49314
rect 1970 49144 2262 49314
rect 2430 49144 2630 49314
rect 2798 49144 3090 49314
rect 3258 49144 3458 49314
rect 3626 49144 3918 49314
rect 4086 49144 4378 49314
rect 4546 49144 4746 49314
rect 4914 49144 5206 49314
rect 5374 49144 5666 49314
rect 5834 49144 6034 49314
rect 6202 49144 6494 49314
rect 6662 49144 6862 49314
rect 7030 49144 7322 49314
rect 7490 49144 7782 49314
rect 7950 49144 8150 49314
rect 8318 49144 8610 49314
rect 8778 49144 8978 49314
rect 9146 49144 9438 49314
rect 9606 49144 9898 49314
rect 10066 49144 10266 49314
rect 10434 49144 10726 49314
rect 10894 49144 11186 49314
rect 11354 49144 11554 49314
rect 11722 49144 12014 49314
rect 12182 49144 12382 49314
rect 12550 49144 12842 49314
rect 13010 49144 13302 49314
rect 13470 49144 13670 49314
rect 13838 49144 14130 49314
rect 14298 49144 14498 49314
rect 14666 49144 14958 49314
rect 15126 49144 15418 49314
rect 15586 49144 15786 49314
rect 15954 49144 16246 49314
rect 16414 49144 16706 49314
rect 16874 49144 17074 49314
rect 17242 49144 17534 49314
rect 17702 49144 17902 49314
rect 18070 49144 18362 49314
rect 18530 49144 18822 49314
rect 18990 49144 19190 49314
rect 19358 49144 19650 49314
rect 20 856 19760 49144
rect 20 800 1342 856
rect 1510 800 4194 856
rect 4362 800 7046 856
rect 7214 800 9898 856
rect 10066 800 12750 856
rect 12918 800 15602 856
rect 15770 800 18454 856
rect 18622 800 19760 856
<< metal3 >>
rect 0 45704 800 45824
rect 19200 43800 20000 43920
rect 0 37408 800 37528
rect 19200 31288 20000 31408
rect 0 29112 800 29232
rect 0 20680 800 20800
rect 19200 18776 20000 18896
rect 0 12384 800 12504
rect 19200 6264 20000 6384
rect 0 4088 800 4208
<< obsm3 >>
rect 800 45904 19200 47361
rect 880 45624 19200 45904
rect 800 44000 19200 45624
rect 800 43720 19120 44000
rect 800 37608 19200 43720
rect 880 37328 19200 37608
rect 800 31488 19200 37328
rect 800 31208 19120 31488
rect 800 29312 19200 31208
rect 880 29032 19200 29312
rect 800 20880 19200 29032
rect 880 20600 19200 20880
rect 800 18976 19200 20600
rect 800 18696 19120 18976
rect 800 12584 19200 18696
rect 880 12304 19200 12584
rect 800 6464 19200 12304
rect 800 6184 19120 6464
rect 800 4288 19200 6184
rect 880 4008 19200 4288
rect 800 2143 19200 4008
<< metal4 >>
rect 3910 2128 4230 47376
rect 6874 2128 7194 47376
rect 9840 2128 10160 47376
rect 12805 2128 13125 47376
rect 15771 2128 16091 47376
<< obsm4 >>
rect 4310 2128 6794 47376
rect 7274 2128 9760 47376
rect 10240 2128 12725 47376
rect 13205 2128 15691 47376
<< labels >>
rlabel metal2 s 14554 49200 14610 50000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 A[2]
port 3 nsew signal input
rlabel metal2 s 16302 49200 16358 50000 6 A[3]
port 4 nsew signal input
rlabel metal2 s 17130 49200 17186 50000 6 A[4]
port 5 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 A[5]
port 6 nsew signal input
rlabel metal3 s 19200 31288 20000 31408 6 A[6]
port 7 nsew signal input
rlabel metal2 s 18418 49200 18474 50000 6 A[7]
port 8 nsew signal input
rlabel metal2 s 18878 49200 18934 50000 6 A[8]
port 9 nsew signal input
rlabel metal2 s 19246 49200 19302 50000 6 A[9]
port 10 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 B[0]
port 11 nsew signal input
rlabel metal3 s 19200 6264 20000 6384 6 B[1]
port 12 nsew signal input
rlabel metal2 s 15474 49200 15530 50000 6 B[2]
port 13 nsew signal input
rlabel metal3 s 19200 18776 20000 18896 6 B[3]
port 14 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 B[4]
port 15 nsew signal input
rlabel metal2 s 17590 49200 17646 50000 6 B[5]
port 16 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 B[6]
port 17 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 B[7]
port 18 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 B[8]
port 19 nsew signal input
rlabel metal2 s 19706 49200 19762 50000 6 B[9]
port 20 nsew signal input
rlabel metal2 s 13726 49200 13782 50000 6 Ci
port 21 nsew signal input
rlabel metal2 s 14186 49200 14242 50000 6 Co
port 22 nsew signal output
rlabel metal2 s 15014 49200 15070 50000 6 S[0]
port 23 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 S[1]
port 24 nsew signal output
rlabel metal2 s 15842 49200 15898 50000 6 S[2]
port 25 nsew signal output
rlabel metal2 s 16762 49200 16818 50000 6 S[3]
port 26 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 S[4]
port 27 nsew signal output
rlabel metal2 s 17958 49200 18014 50000 6 S[5]
port 28 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 S[6]
port 29 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 S[7]
port 30 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 S[8]
port 31 nsew signal output
rlabel metal3 s 19200 43800 20000 43920 6 S[9]
port 32 nsew signal output
rlabel metal2 s 202 49200 258 50000 6 io_oeb[0]
port 33 nsew signal output
rlabel metal2 s 4434 49200 4490 50000 6 io_oeb[10]
port 34 nsew signal output
rlabel metal2 s 4802 49200 4858 50000 6 io_oeb[11]
port 35 nsew signal output
rlabel metal2 s 5262 49200 5318 50000 6 io_oeb[12]
port 36 nsew signal output
rlabel metal2 s 5722 49200 5778 50000 6 io_oeb[13]
port 37 nsew signal output
rlabel metal2 s 6090 49200 6146 50000 6 io_oeb[14]
port 38 nsew signal output
rlabel metal2 s 6550 49200 6606 50000 6 io_oeb[15]
port 39 nsew signal output
rlabel metal2 s 6918 49200 6974 50000 6 io_oeb[16]
port 40 nsew signal output
rlabel metal2 s 7378 49200 7434 50000 6 io_oeb[17]
port 41 nsew signal output
rlabel metal2 s 7838 49200 7894 50000 6 io_oeb[18]
port 42 nsew signal output
rlabel metal2 s 8206 49200 8262 50000 6 io_oeb[19]
port 43 nsew signal output
rlabel metal2 s 570 49200 626 50000 6 io_oeb[1]
port 44 nsew signal output
rlabel metal2 s 8666 49200 8722 50000 6 io_oeb[20]
port 45 nsew signal output
rlabel metal2 s 9034 49200 9090 50000 6 io_oeb[21]
port 46 nsew signal output
rlabel metal2 s 9494 49200 9550 50000 6 io_oeb[22]
port 47 nsew signal output
rlabel metal2 s 9954 49200 10010 50000 6 io_oeb[23]
port 48 nsew signal output
rlabel metal2 s 10322 49200 10378 50000 6 io_oeb[24]
port 49 nsew signal output
rlabel metal2 s 10782 49200 10838 50000 6 io_oeb[25]
port 50 nsew signal output
rlabel metal2 s 11242 49200 11298 50000 6 io_oeb[26]
port 51 nsew signal output
rlabel metal2 s 11610 49200 11666 50000 6 io_oeb[27]
port 52 nsew signal output
rlabel metal2 s 12070 49200 12126 50000 6 io_oeb[28]
port 53 nsew signal output
rlabel metal2 s 12438 49200 12494 50000 6 io_oeb[29]
port 54 nsew signal output
rlabel metal2 s 1030 49200 1086 50000 6 io_oeb[2]
port 55 nsew signal output
rlabel metal2 s 12898 49200 12954 50000 6 io_oeb[30]
port 56 nsew signal output
rlabel metal2 s 13358 49200 13414 50000 6 io_oeb[31]
port 57 nsew signal output
rlabel metal2 s 1398 49200 1454 50000 6 io_oeb[3]
port 58 nsew signal output
rlabel metal2 s 1858 49200 1914 50000 6 io_oeb[4]
port 59 nsew signal output
rlabel metal2 s 2318 49200 2374 50000 6 io_oeb[5]
port 60 nsew signal output
rlabel metal2 s 2686 49200 2742 50000 6 io_oeb[6]
port 61 nsew signal output
rlabel metal2 s 3146 49200 3202 50000 6 io_oeb[7]
port 62 nsew signal output
rlabel metal2 s 3514 49200 3570 50000 6 io_oeb[8]
port 63 nsew signal output
rlabel metal2 s 3974 49200 4030 50000 6 io_oeb[9]
port 64 nsew signal output
rlabel metal4 s 3910 2128 4230 47376 6 vccd1
port 65 nsew power input
rlabel metal4 s 9840 2128 10160 47376 6 vccd1
port 65 nsew power input
rlabel metal4 s 15771 2128 16091 47376 6 vccd1
port 65 nsew power input
rlabel metal4 s 6874 2128 7194 47376 6 vssd1
port 66 nsew ground input
rlabel metal4 s 12805 2128 13125 47376 6 vssd1
port 66 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 813896
string GDS_FILE /home/salah/AI_CORDIC_LIU/mychip/openlane/cordic/runs/cordic/results/finishing/cordic.magic.gds
string GDS_START 200288
<< end >>


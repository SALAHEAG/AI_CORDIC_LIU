magic
tech sky130A
magscale 1 2
timestamp 1695401849
<< viali >>
rect 1501 47209 1535 47243
rect 10241 47209 10275 47243
rect 11529 47209 11563 47243
rect 12173 47209 12207 47243
rect 12817 47209 12851 47243
rect 14657 47141 14691 47175
rect 2145 47073 2179 47107
rect 3801 47073 3835 47107
rect 4445 47073 4479 47107
rect 5089 47073 5123 47107
rect 6377 47073 6411 47107
rect 7665 47073 7699 47107
rect 9597 47073 9631 47107
rect 16129 47073 16163 47107
rect 16681 47073 16715 47107
rect 17969 47073 18003 47107
rect 1685 47005 1719 47039
rect 13553 47005 13587 47039
rect 14841 47005 14875 47039
rect 15853 47005 15887 47039
rect 16957 47005 16991 47039
rect 2789 46937 2823 46971
rect 8953 46937 8987 46971
rect 7021 46869 7055 46903
rect 1409 46665 1443 46699
rect 2053 46665 2087 46699
rect 2697 46665 2731 46699
rect 3525 46665 3559 46699
rect 4905 46665 4939 46699
rect 5549 46665 5583 46699
rect 6745 46665 6779 46699
rect 7665 46665 7699 46699
rect 8585 46665 8619 46699
rect 14197 46665 14231 46699
rect 14933 46665 14967 46699
rect 16681 46665 16715 46699
rect 15761 46597 15795 46631
rect 9505 46529 9539 46563
rect 10517 46529 10551 46563
rect 11897 46529 11931 46563
rect 12817 46529 12851 46563
rect 13461 46529 13495 46563
rect 15117 46529 15151 46563
rect 17601 46529 17635 46563
rect 17325 46461 17359 46495
rect 15577 46393 15611 46427
rect 2053 46121 2087 46155
rect 14105 46121 14139 46155
rect 14749 46121 14783 46155
rect 15485 46121 15519 46155
rect 16313 46121 16347 46155
rect 1409 45985 1443 46019
rect 16957 45985 16991 46019
rect 16497 45917 16531 45951
rect 17233 45917 17267 45951
rect 16129 45509 16163 45543
rect 17141 45441 17175 45475
rect 18061 45441 18095 45475
rect 17325 45305 17359 45339
rect 17877 45305 17911 45339
rect 16865 45033 16899 45067
rect 17417 45033 17451 45067
rect 18061 44829 18095 44863
rect 17877 44761 17911 44795
rect 17969 44489 18003 44523
rect 17417 44421 17451 44455
rect 18153 44353 18187 44387
rect 1685 42177 1719 42211
rect 2145 42177 2179 42211
rect 1501 41973 1535 42007
rect 17509 41089 17543 41123
rect 18153 41089 18187 41123
rect 17969 40885 18003 40919
rect 17969 37213 18003 37247
rect 18153 37213 18187 37247
rect 18061 37145 18095 37179
rect 17049 37077 17083 37111
rect 17141 36873 17175 36907
rect 17969 36805 18003 36839
rect 17325 36737 17359 36771
rect 18153 36737 18187 36771
rect 17785 36533 17819 36567
rect 18061 36329 18095 36363
rect 17693 36193 17727 36227
rect 16681 36125 16715 36159
rect 17785 36125 17819 36159
rect 1869 36057 1903 36091
rect 16497 36057 16531 36091
rect 1961 35989 1995 36023
rect 15669 35989 15703 36023
rect 16313 35989 16347 36023
rect 1685 35785 1719 35819
rect 15485 35785 15519 35819
rect 15301 35649 15335 35683
rect 15945 35649 15979 35683
rect 16129 35649 16163 35683
rect 16681 35649 16715 35683
rect 16865 35649 16899 35683
rect 17693 35649 17727 35683
rect 17785 35581 17819 35615
rect 17325 35513 17359 35547
rect 16037 35445 16071 35479
rect 16773 35445 16807 35479
rect 15209 35105 15243 35139
rect 14381 35037 14415 35071
rect 16589 35037 16623 35071
rect 17417 35037 17451 35071
rect 15945 34969 15979 35003
rect 14289 34697 14323 34731
rect 16865 34697 16899 34731
rect 17417 34629 17451 34663
rect 18061 34629 18095 34663
rect 14105 34561 14139 34595
rect 14289 34561 14323 34595
rect 14749 34561 14783 34595
rect 14933 34561 14967 34595
rect 15761 34561 15795 34595
rect 16681 34561 16715 34595
rect 16957 34561 16991 34595
rect 17785 34561 17819 34595
rect 15669 34493 15703 34527
rect 17877 34493 17911 34527
rect 13645 34425 13679 34459
rect 14841 34425 14875 34459
rect 16129 34425 16163 34459
rect 16681 34357 16715 34391
rect 13461 34153 13495 34187
rect 14473 34153 14507 34187
rect 18061 34153 18095 34187
rect 15853 34085 15887 34119
rect 15577 34017 15611 34051
rect 16405 34017 16439 34051
rect 17325 34017 17359 34051
rect 18153 34017 18187 34051
rect 13369 33949 13403 33983
rect 13553 33949 13587 33983
rect 15485 33949 15519 33983
rect 17233 33949 17267 33983
rect 17877 33949 17911 33983
rect 17969 33949 18003 33983
rect 14657 33881 14691 33915
rect 14841 33881 14875 33915
rect 16497 33881 16531 33915
rect 12725 33813 12759 33847
rect 13829 33609 13863 33643
rect 14289 33541 14323 33575
rect 16129 33541 16163 33575
rect 12725 33473 12759 33507
rect 12817 33473 12851 33507
rect 13461 33473 13495 33507
rect 13645 33473 13679 33507
rect 14473 33473 14507 33507
rect 15491 33473 15525 33507
rect 15648 33479 15682 33513
rect 15761 33473 15795 33507
rect 15853 33473 15887 33507
rect 16957 33473 16991 33507
rect 17417 33473 17451 33507
rect 17785 33473 17819 33507
rect 13001 33405 13035 33439
rect 17509 33405 17543 33439
rect 17417 33337 17451 33371
rect 14657 33269 14691 33303
rect 15117 33065 15151 33099
rect 17233 32929 17267 32963
rect 14289 32861 14323 32895
rect 14381 32861 14415 32895
rect 15301 32861 15335 32895
rect 15393 32861 15427 32895
rect 15485 32861 15519 32895
rect 15577 32861 15611 32895
rect 16313 32861 16347 32895
rect 16497 32861 16531 32895
rect 16865 32861 16899 32895
rect 17325 32861 17359 32895
rect 17693 32861 17727 32895
rect 14565 32793 14599 32827
rect 12909 32725 12943 32759
rect 13461 32725 13495 32759
rect 13645 32521 13679 32555
rect 16129 32521 16163 32555
rect 17417 32521 17451 32555
rect 18061 32521 18095 32555
rect 14105 32385 14139 32419
rect 14289 32385 14323 32419
rect 14749 32385 14783 32419
rect 14841 32385 14875 32419
rect 15025 32385 15059 32419
rect 15669 32385 15703 32419
rect 16681 32385 16715 32419
rect 16865 32385 16899 32419
rect 17141 32385 17175 32419
rect 17877 32385 17911 32419
rect 18061 32385 18095 32419
rect 16957 32249 16991 32283
rect 17049 32249 17083 32283
rect 14105 32181 14139 32215
rect 15209 32181 15243 32215
rect 15945 32181 15979 32215
rect 17233 31977 17267 32011
rect 17601 31909 17635 31943
rect 14749 31841 14783 31875
rect 14105 31773 14139 31807
rect 15669 31773 15703 31807
rect 16405 31773 16439 31807
rect 17141 31773 17175 31807
rect 16681 31433 16715 31467
rect 17969 31433 18003 31467
rect 16037 31365 16071 31399
rect 15393 31297 15427 31331
rect 16865 31297 16899 31331
rect 17049 31297 17083 31331
rect 17141 31297 17175 31331
rect 17601 31297 17635 31331
rect 17693 31297 17727 31331
rect 15209 31229 15243 31263
rect 15577 31161 15611 31195
rect 17601 31093 17635 31127
rect 17417 30889 17451 30923
rect 16865 30821 16899 30855
rect 1409 30685 1443 30719
rect 1685 30685 1719 30719
rect 15853 30685 15887 30719
rect 16037 30685 16071 30719
rect 16589 30685 16623 30719
rect 16681 30685 16715 30719
rect 17325 30685 17359 30719
rect 17509 30685 17543 30719
rect 15945 30549 15979 30583
rect 1409 30345 1443 30379
rect 17325 30345 17359 30379
rect 16773 30277 16807 30311
rect 15761 30209 15795 30243
rect 15853 30209 15887 30243
rect 16681 30209 16715 30243
rect 16865 30209 16899 30243
rect 17325 30209 17359 30243
rect 17509 30209 17543 30243
rect 17969 30209 18003 30243
rect 18153 30209 18187 30243
rect 16037 30073 16071 30107
rect 17969 30073 18003 30107
rect 15853 29597 15887 29631
rect 16037 29597 16071 29631
rect 17785 29597 17819 29631
rect 17969 29597 18003 29631
rect 15945 29529 15979 29563
rect 18061 29461 18095 29495
rect 17969 28713 18003 28747
rect 17509 28509 17543 28543
rect 18153 28509 18187 28543
rect 14381 25993 14415 26027
rect 14105 25857 14139 25891
rect 13737 25789 13771 25823
rect 14197 25789 14231 25823
rect 13185 25449 13219 25483
rect 1685 25245 1719 25279
rect 1501 25109 1535 25143
rect 12817 24837 12851 24871
rect 12633 24769 12667 24803
rect 13461 24769 13495 24803
rect 13645 24769 13679 24803
rect 13001 24701 13035 24735
rect 13553 24565 13587 24599
rect 12633 24361 12667 24395
rect 11161 24293 11195 24327
rect 13185 24293 13219 24327
rect 11621 24225 11655 24259
rect 11529 24157 11563 24191
rect 12541 24157 12575 24191
rect 12725 24157 12759 24191
rect 13553 22049 13587 22083
rect 14105 22049 14139 22083
rect 13277 21981 13311 22015
rect 13369 21981 13403 22015
rect 17509 21981 17543 22015
rect 18153 21981 18187 22015
rect 12909 21845 12943 21879
rect 17969 21845 18003 21879
rect 13277 20417 13311 20451
rect 13461 20417 13495 20451
rect 13369 20213 13403 20247
rect 1685 19873 1719 19907
rect 1409 19805 1443 19839
rect 1409 19397 1443 19431
rect 15301 19329 15335 19363
rect 14473 19261 14507 19295
rect 15209 19261 15243 19295
rect 16129 19261 16163 19295
rect 10977 18377 11011 18411
rect 11897 18377 11931 18411
rect 10333 18241 10367 18275
rect 10793 18241 10827 18275
rect 10977 18241 11011 18275
rect 11529 18241 11563 18275
rect 11713 18241 11747 18275
rect 11345 17493 11379 17527
rect 17877 16065 17911 16099
rect 18153 15997 18187 16031
rect 18153 15657 18187 15691
rect 1685 13889 1719 13923
rect 1409 13821 1443 13855
rect 1409 13481 1443 13515
rect 17417 9537 17451 9571
rect 17877 9537 17911 9571
rect 18061 9401 18095 9435
rect 1869 8449 1903 8483
rect 2053 8313 2087 8347
rect 1593 8041 1627 8075
rect 17877 3485 17911 3519
rect 18061 3349 18095 3383
rect 1685 3009 1719 3043
rect 2237 2941 2271 2975
rect 1501 2805 1535 2839
rect 12725 2601 12759 2635
rect 17693 2601 17727 2635
rect 8401 2533 8435 2567
rect 7849 2397 7883 2431
rect 12081 2397 12115 2431
rect 12541 2397 12575 2431
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 2145 2329 2179 2363
rect 2697 2329 2731 2363
rect 3065 2329 3099 2363
rect 7665 2261 7699 2295
<< metal1 >>
rect 18230 47404 18236 47456
rect 18288 47444 18294 47456
rect 18414 47444 18420 47456
rect 18288 47416 18420 47444
rect 18288 47404 18294 47416
rect 18414 47404 18420 47416
rect 18472 47404 18478 47456
rect 1104 47354 18860 47376
rect 1104 47302 3915 47354
rect 3967 47302 3979 47354
rect 4031 47302 4043 47354
rect 4095 47302 4107 47354
rect 4159 47302 4171 47354
rect 4223 47302 9846 47354
rect 9898 47302 9910 47354
rect 9962 47302 9974 47354
rect 10026 47302 10038 47354
rect 10090 47302 10102 47354
rect 10154 47302 15776 47354
rect 15828 47302 15840 47354
rect 15892 47302 15904 47354
rect 15956 47302 15968 47354
rect 16020 47302 16032 47354
rect 16084 47302 18860 47354
rect 1104 47280 18860 47302
rect 1486 47240 1492 47252
rect 1447 47212 1492 47240
rect 1486 47200 1492 47212
rect 1544 47200 1550 47252
rect 10226 47240 10232 47252
rect 10187 47212 10232 47240
rect 10226 47200 10232 47212
rect 10284 47200 10290 47252
rect 11054 47200 11060 47252
rect 11112 47240 11118 47252
rect 11517 47243 11575 47249
rect 11517 47240 11529 47243
rect 11112 47212 11529 47240
rect 11112 47200 11118 47212
rect 11517 47209 11529 47212
rect 11563 47209 11575 47243
rect 11517 47203 11575 47209
rect 11698 47200 11704 47252
rect 11756 47240 11762 47252
rect 12161 47243 12219 47249
rect 12161 47240 12173 47243
rect 11756 47212 12173 47240
rect 11756 47200 11762 47212
rect 12161 47209 12173 47212
rect 12207 47209 12219 47243
rect 12161 47203 12219 47209
rect 12434 47200 12440 47252
rect 12492 47240 12498 47252
rect 12805 47243 12863 47249
rect 12805 47240 12817 47243
rect 12492 47212 12817 47240
rect 12492 47200 12498 47212
rect 12805 47209 12817 47212
rect 12851 47209 12863 47243
rect 12805 47203 12863 47209
rect 13998 47132 14004 47184
rect 14056 47172 14062 47184
rect 14645 47175 14703 47181
rect 14645 47172 14657 47175
rect 14056 47144 14657 47172
rect 14056 47132 14062 47144
rect 14645 47141 14657 47144
rect 14691 47141 14703 47175
rect 14645 47135 14703 47141
rect 1118 47064 1124 47116
rect 1176 47104 1182 47116
rect 2133 47107 2191 47113
rect 2133 47104 2145 47107
rect 1176 47076 2145 47104
rect 1176 47064 1182 47076
rect 2133 47073 2145 47076
rect 2179 47073 2191 47107
rect 2133 47067 2191 47073
rect 2958 47064 2964 47116
rect 3016 47104 3022 47116
rect 3789 47107 3847 47113
rect 3789 47104 3801 47107
rect 3016 47076 3801 47104
rect 3016 47064 3022 47076
rect 3789 47073 3801 47076
rect 3835 47073 3847 47107
rect 3789 47067 3847 47073
rect 4246 47064 4252 47116
rect 4304 47104 4310 47116
rect 4433 47107 4491 47113
rect 4433 47104 4445 47107
rect 4304 47076 4445 47104
rect 4304 47064 4310 47076
rect 4433 47073 4445 47076
rect 4479 47073 4491 47107
rect 4433 47067 4491 47073
rect 4706 47064 4712 47116
rect 4764 47104 4770 47116
rect 5077 47107 5135 47113
rect 5077 47104 5089 47107
rect 4764 47076 5089 47104
rect 4764 47064 4770 47076
rect 5077 47073 5089 47076
rect 5123 47073 5135 47107
rect 5077 47067 5135 47073
rect 5718 47064 5724 47116
rect 5776 47104 5782 47116
rect 6365 47107 6423 47113
rect 6365 47104 6377 47107
rect 5776 47076 6377 47104
rect 5776 47064 5782 47076
rect 6365 47073 6377 47076
rect 6411 47073 6423 47107
rect 6365 47067 6423 47073
rect 7098 47064 7104 47116
rect 7156 47104 7162 47116
rect 7653 47107 7711 47113
rect 7653 47104 7665 47107
rect 7156 47076 7665 47104
rect 7156 47064 7162 47076
rect 7653 47073 7665 47076
rect 7699 47073 7711 47107
rect 7653 47067 7711 47073
rect 8938 47064 8944 47116
rect 8996 47104 9002 47116
rect 9585 47107 9643 47113
rect 9585 47104 9597 47107
rect 8996 47076 9597 47104
rect 8996 47064 9002 47076
rect 9585 47073 9597 47076
rect 9631 47073 9643 47107
rect 16114 47104 16120 47116
rect 16075 47076 16120 47104
rect 9585 47067 9643 47073
rect 16114 47064 16120 47076
rect 16172 47064 16178 47116
rect 16482 47064 16488 47116
rect 16540 47104 16546 47116
rect 16669 47107 16727 47113
rect 16669 47104 16681 47107
rect 16540 47076 16681 47104
rect 16540 47064 16546 47076
rect 16669 47073 16681 47076
rect 16715 47104 16727 47107
rect 17957 47107 18015 47113
rect 17957 47104 17969 47107
rect 16715 47076 17969 47104
rect 16715 47073 16727 47076
rect 16669 47067 16727 47073
rect 17957 47073 17969 47076
rect 18003 47073 18015 47107
rect 17957 47067 18015 47073
rect 1670 47036 1676 47048
rect 1631 47008 1676 47036
rect 1670 46996 1676 47008
rect 1728 46996 1734 47048
rect 13541 47039 13599 47045
rect 13541 47005 13553 47039
rect 13587 47036 13599 47039
rect 14826 47036 14832 47048
rect 13587 47008 14832 47036
rect 13587 47005 13599 47008
rect 13541 46999 13599 47005
rect 14826 46996 14832 47008
rect 14884 46996 14890 47048
rect 15286 46996 15292 47048
rect 15344 47036 15350 47048
rect 15841 47039 15899 47045
rect 15841 47036 15853 47039
rect 15344 47008 15853 47036
rect 15344 46996 15350 47008
rect 15841 47005 15853 47008
rect 15887 47005 15899 47039
rect 15841 46999 15899 47005
rect 16850 46996 16856 47048
rect 16908 47036 16914 47048
rect 16945 47039 17003 47045
rect 16945 47036 16957 47039
rect 16908 47008 16957 47036
rect 16908 46996 16914 47008
rect 16945 47005 16957 47008
rect 16991 47005 17003 47039
rect 16945 46999 17003 47005
rect 2777 46971 2835 46977
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 2777 46931 2835 46937
rect 8941 46971 8999 46977
rect 8941 46937 8953 46971
rect 8987 46937 8999 46971
rect 8941 46931 8999 46937
rect 2314 46860 2320 46912
rect 2372 46900 2378 46912
rect 2792 46900 2820 46931
rect 2372 46872 2820 46900
rect 2372 46860 2378 46872
rect 6178 46860 6184 46912
rect 6236 46900 6242 46912
rect 7009 46903 7067 46909
rect 7009 46900 7021 46903
rect 6236 46872 7021 46900
rect 6236 46860 6242 46872
rect 7009 46869 7021 46872
rect 7055 46869 7067 46903
rect 7009 46863 7067 46869
rect 8018 46860 8024 46912
rect 8076 46900 8082 46912
rect 8956 46900 8984 46931
rect 8076 46872 8984 46900
rect 8076 46860 8082 46872
rect 1104 46810 18860 46832
rect 1104 46758 6880 46810
rect 6932 46758 6944 46810
rect 6996 46758 7008 46810
rect 7060 46758 7072 46810
rect 7124 46758 7136 46810
rect 7188 46758 12811 46810
rect 12863 46758 12875 46810
rect 12927 46758 12939 46810
rect 12991 46758 13003 46810
rect 13055 46758 13067 46810
rect 13119 46758 18860 46810
rect 1104 46736 18860 46758
rect 658 46656 664 46708
rect 716 46696 722 46708
rect 1397 46699 1455 46705
rect 1397 46696 1409 46699
rect 716 46668 1409 46696
rect 716 46656 722 46668
rect 1397 46665 1409 46668
rect 1443 46665 1455 46699
rect 1397 46659 1455 46665
rect 1578 46656 1584 46708
rect 1636 46696 1642 46708
rect 2041 46699 2099 46705
rect 2041 46696 2053 46699
rect 1636 46668 2053 46696
rect 1636 46656 1642 46668
rect 2041 46665 2053 46668
rect 2087 46665 2099 46699
rect 2682 46696 2688 46708
rect 2643 46668 2688 46696
rect 2041 46659 2099 46665
rect 2682 46656 2688 46668
rect 2740 46656 2746 46708
rect 3510 46696 3516 46708
rect 3471 46668 3516 46696
rect 3510 46656 3516 46668
rect 3568 46656 3574 46708
rect 4890 46696 4896 46708
rect 4851 46668 4896 46696
rect 4890 46656 4896 46668
rect 4948 46656 4954 46708
rect 5258 46656 5264 46708
rect 5316 46696 5322 46708
rect 5537 46699 5595 46705
rect 5537 46696 5549 46699
rect 5316 46668 5549 46696
rect 5316 46656 5322 46668
rect 5537 46665 5549 46668
rect 5583 46665 5595 46699
rect 6730 46696 6736 46708
rect 6691 46668 6736 46696
rect 5537 46659 5595 46665
rect 6730 46656 6736 46668
rect 6788 46656 6794 46708
rect 7650 46696 7656 46708
rect 7611 46668 7656 46696
rect 7650 46656 7656 46668
rect 7708 46656 7714 46708
rect 8570 46696 8576 46708
rect 8531 46668 8576 46696
rect 8570 46656 8576 46668
rect 8628 46656 8634 46708
rect 14182 46696 14188 46708
rect 14143 46668 14188 46696
rect 14182 46656 14188 46668
rect 14240 46656 14246 46708
rect 14921 46699 14979 46705
rect 14921 46665 14933 46699
rect 14967 46696 14979 46699
rect 14967 46668 15884 46696
rect 14967 46665 14979 46668
rect 14921 46659 14979 46665
rect 15470 46588 15476 46640
rect 15528 46628 15534 46640
rect 15749 46631 15807 46637
rect 15749 46628 15761 46631
rect 15528 46600 15761 46628
rect 15528 46588 15534 46600
rect 15749 46597 15761 46600
rect 15795 46597 15807 46631
rect 15856 46628 15884 46668
rect 16114 46656 16120 46708
rect 16172 46696 16178 46708
rect 16669 46699 16727 46705
rect 16669 46696 16681 46699
rect 16172 46668 16681 46696
rect 16172 46656 16178 46668
rect 16669 46665 16681 46668
rect 16715 46665 16727 46699
rect 16669 46659 16727 46665
rect 19150 46628 19156 46640
rect 15856 46600 19156 46628
rect 15749 46591 15807 46597
rect 19150 46588 19156 46600
rect 19208 46588 19214 46640
rect 9490 46560 9496 46572
rect 9451 46532 9496 46560
rect 9490 46520 9496 46532
rect 9548 46520 9554 46572
rect 10502 46560 10508 46572
rect 10463 46532 10508 46560
rect 10502 46520 10508 46532
rect 10560 46520 10566 46572
rect 11882 46560 11888 46572
rect 11843 46532 11888 46560
rect 11882 46520 11888 46532
rect 11940 46520 11946 46572
rect 12710 46520 12716 46572
rect 12768 46560 12774 46572
rect 12805 46563 12863 46569
rect 12805 46560 12817 46563
rect 12768 46532 12817 46560
rect 12768 46520 12774 46532
rect 12805 46529 12817 46532
rect 12851 46529 12863 46563
rect 13446 46560 13452 46572
rect 13407 46532 13452 46560
rect 12805 46523 12863 46529
rect 13446 46520 13452 46532
rect 13504 46520 13510 46572
rect 15102 46560 15108 46572
rect 15063 46532 15108 46560
rect 15102 46520 15108 46532
rect 15160 46520 15166 46572
rect 15654 46520 15660 46572
rect 15712 46560 15718 46572
rect 17589 46563 17647 46569
rect 17589 46560 17601 46563
rect 15712 46532 17601 46560
rect 15712 46520 15718 46532
rect 17589 46529 17601 46532
rect 17635 46529 17647 46563
rect 17589 46523 17647 46529
rect 17310 46492 17316 46504
rect 17223 46464 17316 46492
rect 17310 46452 17316 46464
rect 17368 46492 17374 46504
rect 19610 46492 19616 46504
rect 17368 46464 19616 46492
rect 17368 46452 17374 46464
rect 19610 46452 19616 46464
rect 19668 46452 19674 46504
rect 15562 46424 15568 46436
rect 15523 46396 15568 46424
rect 15562 46384 15568 46396
rect 15620 46384 15626 46436
rect 1104 46266 18860 46288
rect 1104 46214 3915 46266
rect 3967 46214 3979 46266
rect 4031 46214 4043 46266
rect 4095 46214 4107 46266
rect 4159 46214 4171 46266
rect 4223 46214 9846 46266
rect 9898 46214 9910 46266
rect 9962 46214 9974 46266
rect 10026 46214 10038 46266
rect 10090 46214 10102 46266
rect 10154 46214 15776 46266
rect 15828 46214 15840 46266
rect 15892 46214 15904 46266
rect 15956 46214 15968 46266
rect 16020 46214 16032 46266
rect 16084 46214 18860 46266
rect 1104 46192 18860 46214
rect 1670 46112 1676 46164
rect 1728 46152 1734 46164
rect 2038 46152 2044 46164
rect 1728 46124 2044 46152
rect 1728 46112 1734 46124
rect 2038 46112 2044 46124
rect 2096 46112 2102 46164
rect 13630 46112 13636 46164
rect 13688 46152 13694 46164
rect 14093 46155 14151 46161
rect 14093 46152 14105 46155
rect 13688 46124 14105 46152
rect 13688 46112 13694 46124
rect 14093 46121 14105 46124
rect 14139 46121 14151 46155
rect 14734 46152 14740 46164
rect 14695 46124 14740 46152
rect 14093 46115 14151 46121
rect 14734 46112 14740 46124
rect 14792 46112 14798 46164
rect 15470 46152 15476 46164
rect 15431 46124 15476 46152
rect 15470 46112 15476 46124
rect 15528 46112 15534 46164
rect 16301 46155 16359 46161
rect 16301 46121 16313 46155
rect 16347 46152 16359 46155
rect 17770 46152 17776 46164
rect 16347 46124 17776 46152
rect 16347 46121 16359 46124
rect 16301 46115 16359 46121
rect 17770 46112 17776 46124
rect 17828 46112 17834 46164
rect 198 45976 204 46028
rect 256 46016 262 46028
rect 1397 46019 1455 46025
rect 1397 46016 1409 46019
rect 256 45988 1409 46016
rect 256 45976 262 45988
rect 1397 45985 1409 45988
rect 1443 45985 1455 46019
rect 16942 46016 16948 46028
rect 16903 45988 16948 46016
rect 1397 45979 1455 45985
rect 16942 45976 16948 45988
rect 17000 45976 17006 46028
rect 16485 45951 16543 45957
rect 16485 45917 16497 45951
rect 16531 45948 16543 45951
rect 17034 45948 17040 45960
rect 16531 45920 17040 45948
rect 16531 45917 16543 45920
rect 16485 45911 16543 45917
rect 17034 45908 17040 45920
rect 17092 45908 17098 45960
rect 17218 45948 17224 45960
rect 17179 45920 17224 45948
rect 17218 45908 17224 45920
rect 17276 45908 17282 45960
rect 1104 45722 18860 45744
rect 1104 45670 6880 45722
rect 6932 45670 6944 45722
rect 6996 45670 7008 45722
rect 7060 45670 7072 45722
rect 7124 45670 7136 45722
rect 7188 45670 12811 45722
rect 12863 45670 12875 45722
rect 12927 45670 12939 45722
rect 12991 45670 13003 45722
rect 13055 45670 13067 45722
rect 13119 45670 18860 45722
rect 1104 45648 18860 45670
rect 16117 45543 16175 45549
rect 16117 45509 16129 45543
rect 16163 45540 16175 45543
rect 17310 45540 17316 45552
rect 16163 45512 17316 45540
rect 16163 45509 16175 45512
rect 16117 45503 16175 45509
rect 17310 45500 17316 45512
rect 17368 45500 17374 45552
rect 17126 45472 17132 45484
rect 17087 45444 17132 45472
rect 17126 45432 17132 45444
rect 17184 45432 17190 45484
rect 18046 45472 18052 45484
rect 18007 45444 18052 45472
rect 18046 45432 18052 45444
rect 18104 45472 18110 45484
rect 18322 45472 18328 45484
rect 18104 45444 18328 45472
rect 18104 45432 18110 45444
rect 18322 45432 18328 45444
rect 18380 45432 18386 45484
rect 17313 45339 17371 45345
rect 17313 45305 17325 45339
rect 17359 45336 17371 45339
rect 17402 45336 17408 45348
rect 17359 45308 17408 45336
rect 17359 45305 17371 45308
rect 17313 45299 17371 45305
rect 17402 45296 17408 45308
rect 17460 45296 17466 45348
rect 17586 45296 17592 45348
rect 17644 45336 17650 45348
rect 17865 45339 17923 45345
rect 17865 45336 17877 45339
rect 17644 45308 17877 45336
rect 17644 45296 17650 45308
rect 17865 45305 17877 45308
rect 17911 45305 17923 45339
rect 17865 45299 17923 45305
rect 1104 45178 18860 45200
rect 1104 45126 3915 45178
rect 3967 45126 3979 45178
rect 4031 45126 4043 45178
rect 4095 45126 4107 45178
rect 4159 45126 4171 45178
rect 4223 45126 9846 45178
rect 9898 45126 9910 45178
rect 9962 45126 9974 45178
rect 10026 45126 10038 45178
rect 10090 45126 10102 45178
rect 10154 45126 15776 45178
rect 15828 45126 15840 45178
rect 15892 45126 15904 45178
rect 15956 45126 15968 45178
rect 16020 45126 16032 45178
rect 16084 45126 18860 45178
rect 1104 45104 18860 45126
rect 16853 45067 16911 45073
rect 16853 45033 16865 45067
rect 16899 45064 16911 45067
rect 16942 45064 16948 45076
rect 16899 45036 16948 45064
rect 16899 45033 16911 45036
rect 16853 45027 16911 45033
rect 16942 45024 16948 45036
rect 17000 45024 17006 45076
rect 17405 45067 17463 45073
rect 17405 45033 17417 45067
rect 17451 45064 17463 45067
rect 18046 45064 18052 45076
rect 17451 45036 18052 45064
rect 17451 45033 17463 45036
rect 17405 45027 17463 45033
rect 18046 45024 18052 45036
rect 18104 45024 18110 45076
rect 18049 44863 18107 44869
rect 18049 44829 18061 44863
rect 18095 44860 18107 44863
rect 18230 44860 18236 44872
rect 18095 44832 18236 44860
rect 18095 44829 18107 44832
rect 18049 44823 18107 44829
rect 18230 44820 18236 44832
rect 18288 44820 18294 44872
rect 15470 44752 15476 44804
rect 15528 44792 15534 44804
rect 17865 44795 17923 44801
rect 17865 44792 17877 44795
rect 15528 44764 17877 44792
rect 15528 44752 15534 44764
rect 17865 44761 17877 44764
rect 17911 44761 17923 44795
rect 17865 44755 17923 44761
rect 1104 44634 18860 44656
rect 1104 44582 6880 44634
rect 6932 44582 6944 44634
rect 6996 44582 7008 44634
rect 7060 44582 7072 44634
rect 7124 44582 7136 44634
rect 7188 44582 12811 44634
rect 12863 44582 12875 44634
rect 12927 44582 12939 44634
rect 12991 44582 13003 44634
rect 13055 44582 13067 44634
rect 13119 44582 18860 44634
rect 1104 44560 18860 44582
rect 16482 44480 16488 44532
rect 16540 44520 16546 44532
rect 17957 44523 18015 44529
rect 17957 44520 17969 44523
rect 16540 44492 17969 44520
rect 16540 44480 16546 44492
rect 17957 44489 17969 44492
rect 18003 44489 18015 44523
rect 17957 44483 18015 44489
rect 17405 44455 17463 44461
rect 17405 44421 17417 44455
rect 17451 44452 17463 44455
rect 18230 44452 18236 44464
rect 17451 44424 18236 44452
rect 17451 44421 17463 44424
rect 17405 44415 17463 44421
rect 18230 44412 18236 44424
rect 18288 44412 18294 44464
rect 18046 44344 18052 44396
rect 18104 44384 18110 44396
rect 18141 44387 18199 44393
rect 18141 44384 18153 44387
rect 18104 44356 18153 44384
rect 18104 44344 18110 44356
rect 18141 44353 18153 44356
rect 18187 44353 18199 44387
rect 18141 44347 18199 44353
rect 1104 44090 18860 44112
rect 1104 44038 3915 44090
rect 3967 44038 3979 44090
rect 4031 44038 4043 44090
rect 4095 44038 4107 44090
rect 4159 44038 4171 44090
rect 4223 44038 9846 44090
rect 9898 44038 9910 44090
rect 9962 44038 9974 44090
rect 10026 44038 10038 44090
rect 10090 44038 10102 44090
rect 10154 44038 15776 44090
rect 15828 44038 15840 44090
rect 15892 44038 15904 44090
rect 15956 44038 15968 44090
rect 16020 44038 16032 44090
rect 16084 44038 18860 44090
rect 1104 44016 18860 44038
rect 1104 43546 18860 43568
rect 1104 43494 6880 43546
rect 6932 43494 6944 43546
rect 6996 43494 7008 43546
rect 7060 43494 7072 43546
rect 7124 43494 7136 43546
rect 7188 43494 12811 43546
rect 12863 43494 12875 43546
rect 12927 43494 12939 43546
rect 12991 43494 13003 43546
rect 13055 43494 13067 43546
rect 13119 43494 18860 43546
rect 1104 43472 18860 43494
rect 1104 43002 18860 43024
rect 1104 42950 3915 43002
rect 3967 42950 3979 43002
rect 4031 42950 4043 43002
rect 4095 42950 4107 43002
rect 4159 42950 4171 43002
rect 4223 42950 9846 43002
rect 9898 42950 9910 43002
rect 9962 42950 9974 43002
rect 10026 42950 10038 43002
rect 10090 42950 10102 43002
rect 10154 42950 15776 43002
rect 15828 42950 15840 43002
rect 15892 42950 15904 43002
rect 15956 42950 15968 43002
rect 16020 42950 16032 43002
rect 16084 42950 18860 43002
rect 1104 42928 18860 42950
rect 1104 42458 18860 42480
rect 1104 42406 6880 42458
rect 6932 42406 6944 42458
rect 6996 42406 7008 42458
rect 7060 42406 7072 42458
rect 7124 42406 7136 42458
rect 7188 42406 12811 42458
rect 12863 42406 12875 42458
rect 12927 42406 12939 42458
rect 12991 42406 13003 42458
rect 13055 42406 13067 42458
rect 13119 42406 18860 42458
rect 1104 42384 18860 42406
rect 1670 42208 1676 42220
rect 1631 42180 1676 42208
rect 1670 42168 1676 42180
rect 1728 42208 1734 42220
rect 2133 42211 2191 42217
rect 2133 42208 2145 42211
rect 1728 42180 2145 42208
rect 1728 42168 1734 42180
rect 2133 42177 2145 42180
rect 2179 42177 2191 42211
rect 2133 42171 2191 42177
rect 1486 42004 1492 42016
rect 1447 41976 1492 42004
rect 1486 41964 1492 41976
rect 1544 41964 1550 42016
rect 1104 41914 18860 41936
rect 1104 41862 3915 41914
rect 3967 41862 3979 41914
rect 4031 41862 4043 41914
rect 4095 41862 4107 41914
rect 4159 41862 4171 41914
rect 4223 41862 9846 41914
rect 9898 41862 9910 41914
rect 9962 41862 9974 41914
rect 10026 41862 10038 41914
rect 10090 41862 10102 41914
rect 10154 41862 15776 41914
rect 15828 41862 15840 41914
rect 15892 41862 15904 41914
rect 15956 41862 15968 41914
rect 16020 41862 16032 41914
rect 16084 41862 18860 41914
rect 1104 41840 18860 41862
rect 1104 41370 18860 41392
rect 1104 41318 6880 41370
rect 6932 41318 6944 41370
rect 6996 41318 7008 41370
rect 7060 41318 7072 41370
rect 7124 41318 7136 41370
rect 7188 41318 12811 41370
rect 12863 41318 12875 41370
rect 12927 41318 12939 41370
rect 12991 41318 13003 41370
rect 13055 41318 13067 41370
rect 13119 41318 18860 41370
rect 1104 41296 18860 41318
rect 17497 41123 17555 41129
rect 17497 41089 17509 41123
rect 17543 41120 17555 41123
rect 18138 41120 18144 41132
rect 17543 41092 18144 41120
rect 17543 41089 17555 41092
rect 17497 41083 17555 41089
rect 18138 41080 18144 41092
rect 18196 41080 18202 41132
rect 17954 40916 17960 40928
rect 17915 40888 17960 40916
rect 17954 40876 17960 40888
rect 18012 40876 18018 40928
rect 1104 40826 18860 40848
rect 1104 40774 3915 40826
rect 3967 40774 3979 40826
rect 4031 40774 4043 40826
rect 4095 40774 4107 40826
rect 4159 40774 4171 40826
rect 4223 40774 9846 40826
rect 9898 40774 9910 40826
rect 9962 40774 9974 40826
rect 10026 40774 10038 40826
rect 10090 40774 10102 40826
rect 10154 40774 15776 40826
rect 15828 40774 15840 40826
rect 15892 40774 15904 40826
rect 15956 40774 15968 40826
rect 16020 40774 16032 40826
rect 16084 40774 18860 40826
rect 1104 40752 18860 40774
rect 1104 40282 18860 40304
rect 1104 40230 6880 40282
rect 6932 40230 6944 40282
rect 6996 40230 7008 40282
rect 7060 40230 7072 40282
rect 7124 40230 7136 40282
rect 7188 40230 12811 40282
rect 12863 40230 12875 40282
rect 12927 40230 12939 40282
rect 12991 40230 13003 40282
rect 13055 40230 13067 40282
rect 13119 40230 18860 40282
rect 1104 40208 18860 40230
rect 1104 39738 18860 39760
rect 1104 39686 3915 39738
rect 3967 39686 3979 39738
rect 4031 39686 4043 39738
rect 4095 39686 4107 39738
rect 4159 39686 4171 39738
rect 4223 39686 9846 39738
rect 9898 39686 9910 39738
rect 9962 39686 9974 39738
rect 10026 39686 10038 39738
rect 10090 39686 10102 39738
rect 10154 39686 15776 39738
rect 15828 39686 15840 39738
rect 15892 39686 15904 39738
rect 15956 39686 15968 39738
rect 16020 39686 16032 39738
rect 16084 39686 18860 39738
rect 1104 39664 18860 39686
rect 1104 39194 18860 39216
rect 1104 39142 6880 39194
rect 6932 39142 6944 39194
rect 6996 39142 7008 39194
rect 7060 39142 7072 39194
rect 7124 39142 7136 39194
rect 7188 39142 12811 39194
rect 12863 39142 12875 39194
rect 12927 39142 12939 39194
rect 12991 39142 13003 39194
rect 13055 39142 13067 39194
rect 13119 39142 18860 39194
rect 1104 39120 18860 39142
rect 1104 38650 18860 38672
rect 1104 38598 3915 38650
rect 3967 38598 3979 38650
rect 4031 38598 4043 38650
rect 4095 38598 4107 38650
rect 4159 38598 4171 38650
rect 4223 38598 9846 38650
rect 9898 38598 9910 38650
rect 9962 38598 9974 38650
rect 10026 38598 10038 38650
rect 10090 38598 10102 38650
rect 10154 38598 15776 38650
rect 15828 38598 15840 38650
rect 15892 38598 15904 38650
rect 15956 38598 15968 38650
rect 16020 38598 16032 38650
rect 16084 38598 18860 38650
rect 1104 38576 18860 38598
rect 1104 38106 18860 38128
rect 1104 38054 6880 38106
rect 6932 38054 6944 38106
rect 6996 38054 7008 38106
rect 7060 38054 7072 38106
rect 7124 38054 7136 38106
rect 7188 38054 12811 38106
rect 12863 38054 12875 38106
rect 12927 38054 12939 38106
rect 12991 38054 13003 38106
rect 13055 38054 13067 38106
rect 13119 38054 18860 38106
rect 1104 38032 18860 38054
rect 1104 37562 18860 37584
rect 1104 37510 3915 37562
rect 3967 37510 3979 37562
rect 4031 37510 4043 37562
rect 4095 37510 4107 37562
rect 4159 37510 4171 37562
rect 4223 37510 9846 37562
rect 9898 37510 9910 37562
rect 9962 37510 9974 37562
rect 10026 37510 10038 37562
rect 10090 37510 10102 37562
rect 10154 37510 15776 37562
rect 15828 37510 15840 37562
rect 15892 37510 15904 37562
rect 15956 37510 15968 37562
rect 16020 37510 16032 37562
rect 16084 37510 18860 37562
rect 1104 37488 18860 37510
rect 17954 37244 17960 37256
rect 17915 37216 17960 37244
rect 17954 37204 17960 37216
rect 18012 37204 18018 37256
rect 18138 37244 18144 37256
rect 18099 37216 18144 37244
rect 18138 37204 18144 37216
rect 18196 37204 18202 37256
rect 16390 37136 16396 37188
rect 16448 37176 16454 37188
rect 18049 37179 18107 37185
rect 18049 37176 18061 37179
rect 16448 37148 18061 37176
rect 16448 37136 16454 37148
rect 18049 37145 18061 37148
rect 18095 37145 18107 37179
rect 18049 37139 18107 37145
rect 16942 37068 16948 37120
rect 17000 37108 17006 37120
rect 17037 37111 17095 37117
rect 17037 37108 17049 37111
rect 17000 37080 17049 37108
rect 17000 37068 17006 37080
rect 17037 37077 17049 37080
rect 17083 37077 17095 37111
rect 17037 37071 17095 37077
rect 1104 37018 18860 37040
rect 1104 36966 6880 37018
rect 6932 36966 6944 37018
rect 6996 36966 7008 37018
rect 7060 36966 7072 37018
rect 7124 36966 7136 37018
rect 7188 36966 12811 37018
rect 12863 36966 12875 37018
rect 12927 36966 12939 37018
rect 12991 36966 13003 37018
rect 13055 36966 13067 37018
rect 13119 36966 18860 37018
rect 1104 36944 18860 36966
rect 17034 36864 17040 36916
rect 17092 36904 17098 36916
rect 17129 36907 17187 36913
rect 17129 36904 17141 36907
rect 17092 36876 17141 36904
rect 17092 36864 17098 36876
rect 17129 36873 17141 36876
rect 17175 36873 17187 36907
rect 17129 36867 17187 36873
rect 17954 36836 17960 36848
rect 17915 36808 17960 36836
rect 17954 36796 17960 36808
rect 18012 36796 18018 36848
rect 17313 36771 17371 36777
rect 17313 36737 17325 36771
rect 17359 36737 17371 36771
rect 18138 36768 18144 36780
rect 18099 36740 18144 36768
rect 17313 36731 17371 36737
rect 17328 36700 17356 36731
rect 18138 36728 18144 36740
rect 18196 36728 18202 36780
rect 18230 36700 18236 36712
rect 17328 36672 18236 36700
rect 18230 36660 18236 36672
rect 18288 36660 18294 36712
rect 17770 36564 17776 36576
rect 17731 36536 17776 36564
rect 17770 36524 17776 36536
rect 17828 36524 17834 36576
rect 1104 36474 18860 36496
rect 1104 36422 3915 36474
rect 3967 36422 3979 36474
rect 4031 36422 4043 36474
rect 4095 36422 4107 36474
rect 4159 36422 4171 36474
rect 4223 36422 9846 36474
rect 9898 36422 9910 36474
rect 9962 36422 9974 36474
rect 10026 36422 10038 36474
rect 10090 36422 10102 36474
rect 10154 36422 15776 36474
rect 15828 36422 15840 36474
rect 15892 36422 15904 36474
rect 15956 36422 15968 36474
rect 16020 36422 16032 36474
rect 16084 36422 18860 36474
rect 1104 36400 18860 36422
rect 18046 36360 18052 36372
rect 18007 36332 18052 36360
rect 18046 36320 18052 36332
rect 18104 36320 18110 36372
rect 15194 36184 15200 36236
rect 15252 36224 15258 36236
rect 17681 36227 17739 36233
rect 17681 36224 17693 36227
rect 15252 36196 17693 36224
rect 15252 36184 15258 36196
rect 17681 36193 17693 36196
rect 17727 36193 17739 36227
rect 17681 36187 17739 36193
rect 16669 36159 16727 36165
rect 16669 36125 16681 36159
rect 16715 36156 16727 36159
rect 16850 36156 16856 36168
rect 16715 36128 16856 36156
rect 16715 36125 16727 36128
rect 16669 36119 16727 36125
rect 16850 36116 16856 36128
rect 16908 36116 16914 36168
rect 17773 36159 17831 36165
rect 17773 36125 17785 36159
rect 17819 36156 17831 36159
rect 17954 36156 17960 36168
rect 17819 36128 17960 36156
rect 17819 36125 17831 36128
rect 17773 36119 17831 36125
rect 17954 36116 17960 36128
rect 18012 36116 18018 36168
rect 1854 36088 1860 36100
rect 1815 36060 1860 36088
rect 1854 36048 1860 36060
rect 1912 36048 1918 36100
rect 16485 36091 16543 36097
rect 16485 36057 16497 36091
rect 16531 36088 16543 36091
rect 16574 36088 16580 36100
rect 16531 36060 16580 36088
rect 16531 36057 16543 36060
rect 16485 36051 16543 36057
rect 16574 36048 16580 36060
rect 16632 36088 16638 36100
rect 17218 36088 17224 36100
rect 16632 36060 17224 36088
rect 16632 36048 16638 36060
rect 17218 36048 17224 36060
rect 17276 36048 17282 36100
rect 1949 36023 2007 36029
rect 1949 35989 1961 36023
rect 1995 36020 2007 36023
rect 14274 36020 14280 36032
rect 1995 35992 14280 36020
rect 1995 35989 2007 35992
rect 1949 35983 2007 35989
rect 14274 35980 14280 35992
rect 14332 35980 14338 36032
rect 15654 36020 15660 36032
rect 15615 35992 15660 36020
rect 15654 35980 15660 35992
rect 15712 35980 15718 36032
rect 16298 36020 16304 36032
rect 16259 35992 16304 36020
rect 16298 35980 16304 35992
rect 16356 35980 16362 36032
rect 1104 35930 18860 35952
rect 1104 35878 6880 35930
rect 6932 35878 6944 35930
rect 6996 35878 7008 35930
rect 7060 35878 7072 35930
rect 7124 35878 7136 35930
rect 7188 35878 12811 35930
rect 12863 35878 12875 35930
rect 12927 35878 12939 35930
rect 12991 35878 13003 35930
rect 13055 35878 13067 35930
rect 13119 35878 18860 35930
rect 1104 35856 18860 35878
rect 1673 35819 1731 35825
rect 1673 35785 1685 35819
rect 1719 35816 1731 35819
rect 1854 35816 1860 35828
rect 1719 35788 1860 35816
rect 1719 35785 1731 35788
rect 1673 35779 1731 35785
rect 1854 35776 1860 35788
rect 1912 35776 1918 35828
rect 15473 35819 15531 35825
rect 15473 35785 15485 35819
rect 15519 35816 15531 35819
rect 18138 35816 18144 35828
rect 15519 35788 18144 35816
rect 15519 35785 15531 35788
rect 15473 35779 15531 35785
rect 18138 35776 18144 35788
rect 18196 35776 18202 35828
rect 15562 35708 15568 35760
rect 15620 35748 15626 35760
rect 15620 35720 16160 35748
rect 15620 35708 15626 35720
rect 15289 35683 15347 35689
rect 15289 35649 15301 35683
rect 15335 35680 15347 35683
rect 15654 35680 15660 35692
rect 15335 35652 15660 35680
rect 15335 35649 15347 35652
rect 15289 35643 15347 35649
rect 15654 35640 15660 35652
rect 15712 35640 15718 35692
rect 16132 35689 16160 35720
rect 15933 35683 15991 35689
rect 15933 35649 15945 35683
rect 15979 35649 15991 35683
rect 15933 35643 15991 35649
rect 16117 35683 16175 35689
rect 16117 35649 16129 35683
rect 16163 35649 16175 35683
rect 16117 35643 16175 35649
rect 15948 35612 15976 35643
rect 16574 35640 16580 35692
rect 16632 35680 16638 35692
rect 16669 35683 16727 35689
rect 16669 35680 16681 35683
rect 16632 35652 16681 35680
rect 16632 35640 16638 35652
rect 16669 35649 16681 35652
rect 16715 35649 16727 35683
rect 16850 35680 16856 35692
rect 16811 35652 16856 35680
rect 16669 35643 16727 35649
rect 16850 35640 16856 35652
rect 16908 35640 16914 35692
rect 17034 35640 17040 35692
rect 17092 35680 17098 35692
rect 17681 35683 17739 35689
rect 17681 35680 17693 35683
rect 17092 35652 17693 35680
rect 17092 35640 17098 35652
rect 17681 35649 17693 35652
rect 17727 35649 17739 35683
rect 17681 35643 17739 35649
rect 16206 35612 16212 35624
rect 15948 35584 16212 35612
rect 16206 35572 16212 35584
rect 16264 35572 16270 35624
rect 17773 35615 17831 35621
rect 17773 35581 17785 35615
rect 17819 35612 17831 35615
rect 18046 35612 18052 35624
rect 17819 35584 18052 35612
rect 17819 35581 17831 35584
rect 17773 35575 17831 35581
rect 18046 35572 18052 35584
rect 18104 35572 18110 35624
rect 15102 35504 15108 35556
rect 15160 35544 15166 35556
rect 17313 35547 17371 35553
rect 17313 35544 17325 35547
rect 15160 35516 17325 35544
rect 15160 35504 15166 35516
rect 17313 35513 17325 35516
rect 17359 35513 17371 35547
rect 17313 35507 17371 35513
rect 14458 35436 14464 35488
rect 14516 35476 14522 35488
rect 16025 35479 16083 35485
rect 16025 35476 16037 35479
rect 14516 35448 16037 35476
rect 14516 35436 14522 35448
rect 16025 35445 16037 35448
rect 16071 35445 16083 35479
rect 16025 35439 16083 35445
rect 16761 35479 16819 35485
rect 16761 35445 16773 35479
rect 16807 35476 16819 35479
rect 16850 35476 16856 35488
rect 16807 35448 16856 35476
rect 16807 35445 16819 35448
rect 16761 35439 16819 35445
rect 16850 35436 16856 35448
rect 16908 35436 16914 35488
rect 1104 35386 18860 35408
rect 1104 35334 3915 35386
rect 3967 35334 3979 35386
rect 4031 35334 4043 35386
rect 4095 35334 4107 35386
rect 4159 35334 4171 35386
rect 4223 35334 9846 35386
rect 9898 35334 9910 35386
rect 9962 35334 9974 35386
rect 10026 35334 10038 35386
rect 10090 35334 10102 35386
rect 10154 35334 15776 35386
rect 15828 35334 15840 35386
rect 15892 35334 15904 35386
rect 15956 35334 15968 35386
rect 16020 35334 16032 35386
rect 16084 35334 18860 35386
rect 1104 35312 18860 35334
rect 17494 35272 17500 35284
rect 16408 35244 17500 35272
rect 14366 35164 14372 35216
rect 14424 35204 14430 35216
rect 16022 35204 16028 35216
rect 14424 35176 16028 35204
rect 14424 35164 14430 35176
rect 16022 35164 16028 35176
rect 16080 35164 16086 35216
rect 14826 35096 14832 35148
rect 14884 35136 14890 35148
rect 15197 35139 15255 35145
rect 15197 35136 15209 35139
rect 14884 35108 15209 35136
rect 14884 35096 14890 35108
rect 15197 35105 15209 35108
rect 15243 35136 15255 35139
rect 16408 35136 16436 35244
rect 17494 35232 17500 35244
rect 17552 35232 17558 35284
rect 15243 35108 16436 35136
rect 15243 35105 15255 35108
rect 15197 35099 15255 35105
rect 1670 35028 1676 35080
rect 1728 35068 1734 35080
rect 14369 35071 14427 35077
rect 14369 35068 14381 35071
rect 1728 35040 14381 35068
rect 1728 35028 1734 35040
rect 14369 35037 14381 35040
rect 14415 35037 14427 35071
rect 14369 35031 14427 35037
rect 15102 35028 15108 35080
rect 15160 35028 15166 35080
rect 16574 35068 16580 35080
rect 15856 35040 16436 35068
rect 16535 35040 16580 35068
rect 2038 34960 2044 35012
rect 2096 35000 2102 35012
rect 2096 34972 6914 35000
rect 2096 34960 2102 34972
rect 6886 34932 6914 34972
rect 14918 34960 14924 35012
rect 14976 35000 14982 35012
rect 15856 35000 15884 35040
rect 14976 34972 15884 35000
rect 15933 35003 15991 35009
rect 14976 34960 14982 34972
rect 15933 34969 15945 35003
rect 15979 34969 15991 35003
rect 16408 35000 16436 35040
rect 16574 35028 16580 35040
rect 16632 35028 16638 35080
rect 17405 35071 17463 35077
rect 17405 35037 17417 35071
rect 17451 35068 17463 35071
rect 17862 35068 17868 35080
rect 17451 35040 17868 35068
rect 17451 35037 17463 35040
rect 17405 35031 17463 35037
rect 17862 35028 17868 35040
rect 17920 35028 17926 35080
rect 18138 35000 18144 35012
rect 16408 34972 18144 35000
rect 15933 34963 15991 34969
rect 15948 34932 15976 34963
rect 18138 34960 18144 34972
rect 18196 34960 18202 35012
rect 6886 34904 15976 34932
rect 16022 34892 16028 34944
rect 16080 34932 16086 34944
rect 17770 34932 17776 34944
rect 16080 34904 17776 34932
rect 16080 34892 16086 34904
rect 17770 34892 17776 34904
rect 17828 34892 17834 34944
rect 1104 34842 18860 34864
rect 1104 34790 6880 34842
rect 6932 34790 6944 34842
rect 6996 34790 7008 34842
rect 7060 34790 7072 34842
rect 7124 34790 7136 34842
rect 7188 34790 12811 34842
rect 12863 34790 12875 34842
rect 12927 34790 12939 34842
rect 12991 34790 13003 34842
rect 13055 34790 13067 34842
rect 13119 34790 18860 34842
rect 1104 34768 18860 34790
rect 14277 34731 14335 34737
rect 14277 34697 14289 34731
rect 14323 34728 14335 34731
rect 15194 34728 15200 34740
rect 14323 34700 15200 34728
rect 14323 34697 14335 34700
rect 14277 34691 14335 34697
rect 15194 34688 15200 34700
rect 15252 34688 15258 34740
rect 15470 34688 15476 34740
rect 15528 34728 15534 34740
rect 16853 34731 16911 34737
rect 16853 34728 16865 34731
rect 15528 34700 16865 34728
rect 15528 34688 15534 34700
rect 16853 34697 16865 34700
rect 16899 34697 16911 34731
rect 16853 34691 16911 34697
rect 14458 34620 14464 34672
rect 14516 34660 14522 34672
rect 17405 34663 17463 34669
rect 17405 34660 17417 34663
rect 14516 34632 17417 34660
rect 14516 34620 14522 34632
rect 17405 34629 17417 34632
rect 17451 34629 17463 34663
rect 17405 34623 17463 34629
rect 17954 34620 17960 34672
rect 18012 34660 18018 34672
rect 18049 34663 18107 34669
rect 18049 34660 18061 34663
rect 18012 34632 18061 34660
rect 18012 34620 18018 34632
rect 18049 34629 18061 34632
rect 18095 34629 18107 34663
rect 18049 34623 18107 34629
rect 14093 34595 14151 34601
rect 14093 34561 14105 34595
rect 14139 34561 14151 34595
rect 14093 34555 14151 34561
rect 14277 34595 14335 34601
rect 14277 34561 14289 34595
rect 14323 34592 14335 34595
rect 14366 34592 14372 34604
rect 14323 34564 14372 34592
rect 14323 34561 14335 34564
rect 14277 34555 14335 34561
rect 14108 34524 14136 34555
rect 14366 34552 14372 34564
rect 14424 34552 14430 34604
rect 14734 34592 14740 34604
rect 14695 34564 14740 34592
rect 14734 34552 14740 34564
rect 14792 34552 14798 34604
rect 14918 34592 14924 34604
rect 14879 34564 14924 34592
rect 14918 34552 14924 34564
rect 14976 34552 14982 34604
rect 15010 34552 15016 34604
rect 15068 34592 15074 34604
rect 15749 34595 15807 34601
rect 15749 34592 15761 34595
rect 15068 34564 15761 34592
rect 15068 34552 15074 34564
rect 15749 34561 15761 34564
rect 15795 34561 15807 34595
rect 16390 34592 16396 34604
rect 15749 34555 15807 34561
rect 15856 34564 16396 34592
rect 14108 34496 15240 34524
rect 13630 34456 13636 34468
rect 13591 34428 13636 34456
rect 13630 34416 13636 34428
rect 13688 34416 13694 34468
rect 14826 34456 14832 34468
rect 14787 34428 14832 34456
rect 14826 34416 14832 34428
rect 14884 34416 14890 34468
rect 15212 34456 15240 34496
rect 15378 34484 15384 34536
rect 15436 34524 15442 34536
rect 15657 34527 15715 34533
rect 15657 34524 15669 34527
rect 15436 34496 15669 34524
rect 15436 34484 15442 34496
rect 15657 34493 15669 34496
rect 15703 34493 15715 34527
rect 15657 34487 15715 34493
rect 15856 34456 15884 34564
rect 16390 34552 16396 34564
rect 16448 34552 16454 34604
rect 16669 34595 16727 34601
rect 16669 34561 16681 34595
rect 16715 34592 16727 34595
rect 16758 34592 16764 34604
rect 16715 34564 16764 34592
rect 16715 34561 16727 34564
rect 16669 34555 16727 34561
rect 16758 34552 16764 34564
rect 16816 34552 16822 34604
rect 16942 34592 16948 34604
rect 16903 34564 16948 34592
rect 16942 34552 16948 34564
rect 17000 34552 17006 34604
rect 17773 34595 17831 34601
rect 17773 34561 17785 34595
rect 17819 34561 17831 34595
rect 17773 34555 17831 34561
rect 16482 34484 16488 34536
rect 16540 34524 16546 34536
rect 17788 34524 17816 34555
rect 16540 34496 17816 34524
rect 16540 34484 16546 34496
rect 17862 34484 17868 34536
rect 17920 34524 17926 34536
rect 17920 34496 17965 34524
rect 17920 34484 17926 34496
rect 15212 34428 15884 34456
rect 16117 34459 16175 34465
rect 16117 34425 16129 34459
rect 16163 34456 16175 34459
rect 17126 34456 17132 34468
rect 16163 34428 17132 34456
rect 16163 34425 16175 34428
rect 16117 34419 16175 34425
rect 17126 34416 17132 34428
rect 17184 34416 17190 34468
rect 13446 34348 13452 34400
rect 13504 34388 13510 34400
rect 16574 34388 16580 34400
rect 13504 34360 16580 34388
rect 13504 34348 13510 34360
rect 16574 34348 16580 34360
rect 16632 34348 16638 34400
rect 16669 34391 16727 34397
rect 16669 34357 16681 34391
rect 16715 34388 16727 34391
rect 16942 34388 16948 34400
rect 16715 34360 16948 34388
rect 16715 34357 16727 34360
rect 16669 34351 16727 34357
rect 16942 34348 16948 34360
rect 17000 34348 17006 34400
rect 1104 34298 18860 34320
rect 1104 34246 3915 34298
rect 3967 34246 3979 34298
rect 4031 34246 4043 34298
rect 4095 34246 4107 34298
rect 4159 34246 4171 34298
rect 4223 34246 9846 34298
rect 9898 34246 9910 34298
rect 9962 34246 9974 34298
rect 10026 34246 10038 34298
rect 10090 34246 10102 34298
rect 10154 34246 15776 34298
rect 15828 34246 15840 34298
rect 15892 34246 15904 34298
rect 15956 34246 15968 34298
rect 16020 34246 16032 34298
rect 16084 34246 18860 34298
rect 1104 34224 18860 34246
rect 13446 34184 13452 34196
rect 13407 34156 13452 34184
rect 13446 34144 13452 34156
rect 13504 34144 13510 34196
rect 14461 34187 14519 34193
rect 14461 34153 14473 34187
rect 14507 34184 14519 34187
rect 16482 34184 16488 34196
rect 14507 34156 16488 34184
rect 14507 34153 14519 34156
rect 14461 34147 14519 34153
rect 14476 34116 14504 34147
rect 16482 34144 16488 34156
rect 16540 34144 16546 34196
rect 18046 34184 18052 34196
rect 18007 34156 18052 34184
rect 18046 34144 18052 34156
rect 18104 34144 18110 34196
rect 13372 34088 14504 34116
rect 15841 34119 15899 34125
rect 13372 33989 13400 34088
rect 15841 34085 15853 34119
rect 15887 34085 15899 34119
rect 17954 34116 17960 34128
rect 15841 34079 15899 34085
rect 17328 34088 17960 34116
rect 13630 34008 13636 34060
rect 13688 34048 13694 34060
rect 15565 34051 15623 34057
rect 15565 34048 15577 34051
rect 13688 34020 15577 34048
rect 13688 34008 13694 34020
rect 15565 34017 15577 34020
rect 15611 34048 15623 34051
rect 15654 34048 15660 34060
rect 15611 34020 15660 34048
rect 15611 34017 15623 34020
rect 15565 34011 15623 34017
rect 15654 34008 15660 34020
rect 15712 34048 15718 34060
rect 15856 34048 15884 34079
rect 16390 34048 16396 34060
rect 15712 34020 15792 34048
rect 15856 34020 16252 34048
rect 16351 34020 16396 34048
rect 15712 34008 15718 34020
rect 13357 33983 13415 33989
rect 13357 33949 13369 33983
rect 13403 33949 13415 33983
rect 13357 33943 13415 33949
rect 13541 33983 13599 33989
rect 13541 33949 13553 33983
rect 13587 33980 13599 33983
rect 14458 33980 14464 33992
rect 13587 33952 14464 33980
rect 13587 33949 13599 33952
rect 13541 33943 13599 33949
rect 14458 33940 14464 33952
rect 14516 33940 14522 33992
rect 15470 33980 15476 33992
rect 15431 33952 15476 33980
rect 15470 33940 15476 33952
rect 15528 33940 15534 33992
rect 15764 33980 15792 34020
rect 16022 33980 16028 33992
rect 15764 33952 16028 33980
rect 16022 33940 16028 33952
rect 16080 33940 16086 33992
rect 16224 33980 16252 34020
rect 16390 34008 16396 34020
rect 16448 34008 16454 34060
rect 17328 34057 17356 34088
rect 17954 34076 17960 34088
rect 18012 34076 18018 34128
rect 17313 34051 17371 34057
rect 17313 34017 17325 34051
rect 17359 34017 17371 34051
rect 17313 34011 17371 34017
rect 17494 34008 17500 34060
rect 17552 34048 17558 34060
rect 17678 34048 17684 34060
rect 17552 34020 17684 34048
rect 17552 34008 17558 34020
rect 17678 34008 17684 34020
rect 17736 34048 17742 34060
rect 18138 34048 18144 34060
rect 17736 34020 17908 34048
rect 18099 34020 18144 34048
rect 17736 34008 17742 34020
rect 16666 33980 16672 33992
rect 16224 33952 16672 33980
rect 16666 33940 16672 33952
rect 16724 33980 16730 33992
rect 17034 33980 17040 33992
rect 16724 33952 17040 33980
rect 16724 33940 16730 33952
rect 17034 33940 17040 33952
rect 17092 33940 17098 33992
rect 17221 33983 17279 33989
rect 17221 33949 17233 33983
rect 17267 33980 17279 33983
rect 17770 33980 17776 33992
rect 17267 33952 17776 33980
rect 17267 33949 17279 33952
rect 17221 33943 17279 33949
rect 17770 33940 17776 33952
rect 17828 33940 17834 33992
rect 17880 33989 17908 34020
rect 18138 34008 18144 34020
rect 18196 34008 18202 34060
rect 17865 33983 17923 33989
rect 17865 33949 17877 33983
rect 17911 33949 17923 33983
rect 17865 33943 17923 33949
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33949 18015 33983
rect 17957 33943 18015 33949
rect 14642 33872 14648 33924
rect 14700 33912 14706 33924
rect 14829 33915 14887 33921
rect 14700 33884 14745 33912
rect 14700 33872 14706 33884
rect 14829 33881 14841 33915
rect 14875 33912 14887 33915
rect 15562 33912 15568 33924
rect 14875 33884 15568 33912
rect 14875 33881 14887 33884
rect 14829 33875 14887 33881
rect 15562 33872 15568 33884
rect 15620 33872 15626 33924
rect 16485 33915 16543 33921
rect 15764 33884 16436 33912
rect 12710 33844 12716 33856
rect 12671 33816 12716 33844
rect 12710 33804 12716 33816
rect 12768 33844 12774 33856
rect 13446 33844 13452 33856
rect 12768 33816 13452 33844
rect 12768 33804 12774 33816
rect 13446 33804 13452 33816
rect 13504 33844 13510 33856
rect 14918 33844 14924 33856
rect 13504 33816 14924 33844
rect 13504 33804 13510 33816
rect 14918 33804 14924 33816
rect 14976 33804 14982 33856
rect 15102 33804 15108 33856
rect 15160 33844 15166 33856
rect 15764 33844 15792 33884
rect 15160 33816 15792 33844
rect 16408 33844 16436 33884
rect 16485 33881 16497 33915
rect 16531 33912 16543 33915
rect 16574 33912 16580 33924
rect 16531 33884 16580 33912
rect 16531 33881 16543 33884
rect 16485 33875 16543 33881
rect 16574 33872 16580 33884
rect 16632 33872 16638 33924
rect 17972 33844 18000 33943
rect 16408 33816 18000 33844
rect 15160 33804 15166 33816
rect 1104 33754 18860 33776
rect 1104 33702 6880 33754
rect 6932 33702 6944 33754
rect 6996 33702 7008 33754
rect 7060 33702 7072 33754
rect 7124 33702 7136 33754
rect 7188 33702 12811 33754
rect 12863 33702 12875 33754
rect 12927 33702 12939 33754
rect 12991 33702 13003 33754
rect 13055 33702 13067 33754
rect 13119 33702 18860 33754
rect 1104 33680 18860 33702
rect 13817 33643 13875 33649
rect 13817 33609 13829 33643
rect 13863 33640 13875 33643
rect 14734 33640 14740 33652
rect 13863 33612 14740 33640
rect 13863 33609 13875 33612
rect 13817 33603 13875 33609
rect 14734 33600 14740 33612
rect 14792 33600 14798 33652
rect 14918 33600 14924 33652
rect 14976 33640 14982 33652
rect 14976 33612 15332 33640
rect 14976 33600 14982 33612
rect 14274 33572 14280 33584
rect 12728 33544 13768 33572
rect 14235 33544 14280 33572
rect 12728 33513 12756 33544
rect 12713 33507 12771 33513
rect 12713 33473 12725 33507
rect 12759 33473 12771 33507
rect 12713 33467 12771 33473
rect 12805 33507 12863 33513
rect 12805 33473 12817 33507
rect 12851 33504 12863 33507
rect 13446 33504 13452 33516
rect 12851 33476 12940 33504
rect 13407 33476 13452 33504
rect 12851 33473 12863 33476
rect 12805 33467 12863 33473
rect 12912 33368 12940 33476
rect 13446 33464 13452 33476
rect 13504 33464 13510 33516
rect 13538 33464 13544 33516
rect 13596 33504 13602 33516
rect 13633 33507 13691 33513
rect 13633 33504 13645 33507
rect 13596 33476 13645 33504
rect 13596 33464 13602 33476
rect 13633 33473 13645 33476
rect 13679 33473 13691 33507
rect 13740 33504 13768 33544
rect 14274 33532 14280 33544
rect 14332 33532 14338 33584
rect 15194 33572 15200 33584
rect 14384 33544 15200 33572
rect 14384 33504 14412 33544
rect 15194 33532 15200 33544
rect 15252 33532 15258 33584
rect 13740 33476 14412 33504
rect 14461 33507 14519 33513
rect 13633 33467 13691 33473
rect 14461 33473 14473 33507
rect 14507 33504 14519 33507
rect 14550 33504 14556 33516
rect 14507 33476 14556 33504
rect 14507 33473 14519 33476
rect 14461 33467 14519 33473
rect 14550 33464 14556 33476
rect 14608 33464 14614 33516
rect 14642 33464 14648 33516
rect 14700 33504 14706 33516
rect 15304 33504 15332 33612
rect 15562 33600 15568 33652
rect 15620 33600 15626 33652
rect 15479 33507 15537 33513
rect 15479 33504 15491 33507
rect 14700 33476 15148 33504
rect 15304 33476 15491 33504
rect 14700 33464 14706 33476
rect 12989 33439 13047 33445
rect 12989 33405 13001 33439
rect 13035 33436 13047 33439
rect 15010 33436 15016 33448
rect 13035 33408 15016 33436
rect 13035 33405 13047 33408
rect 12989 33399 13047 33405
rect 15010 33396 15016 33408
rect 15068 33396 15074 33448
rect 15120 33436 15148 33476
rect 15479 33473 15491 33476
rect 15525 33473 15537 33507
rect 15580 33510 15608 33600
rect 16022 33572 16028 33584
rect 15764 33544 16028 33572
rect 15636 33513 15694 33519
rect 15764 33513 15792 33544
rect 16022 33532 16028 33544
rect 16080 33532 16086 33584
rect 16117 33575 16175 33581
rect 16117 33541 16129 33575
rect 16163 33572 16175 33575
rect 16758 33572 16764 33584
rect 16163 33544 16764 33572
rect 16163 33541 16175 33544
rect 16117 33535 16175 33541
rect 16758 33532 16764 33544
rect 16816 33532 16822 33584
rect 15636 33510 15648 33513
rect 15580 33482 15648 33510
rect 15636 33479 15648 33482
rect 15682 33479 15694 33513
rect 15636 33473 15694 33479
rect 15749 33507 15807 33513
rect 15749 33473 15761 33507
rect 15795 33473 15807 33507
rect 15479 33467 15537 33473
rect 15749 33467 15807 33473
rect 15838 33464 15844 33516
rect 15896 33504 15902 33516
rect 16942 33504 16948 33516
rect 15896 33476 15941 33504
rect 16903 33476 16948 33504
rect 15896 33464 15902 33476
rect 16942 33464 16948 33476
rect 17000 33464 17006 33516
rect 17402 33504 17408 33516
rect 17363 33476 17408 33504
rect 17402 33464 17408 33476
rect 17460 33464 17466 33516
rect 17773 33507 17831 33513
rect 17773 33473 17785 33507
rect 17819 33504 17831 33507
rect 17954 33504 17960 33516
rect 17819 33476 17960 33504
rect 17819 33473 17831 33476
rect 17773 33467 17831 33473
rect 17954 33464 17960 33476
rect 18012 33464 18018 33516
rect 16206 33436 16212 33448
rect 15120 33408 16212 33436
rect 16206 33396 16212 33408
rect 16264 33396 16270 33448
rect 17494 33436 17500 33448
rect 17455 33408 17500 33436
rect 17494 33396 17500 33408
rect 17552 33396 17558 33448
rect 16850 33368 16856 33380
rect 12912 33340 16856 33368
rect 16850 33328 16856 33340
rect 16908 33328 16914 33380
rect 17405 33371 17463 33377
rect 17405 33337 17417 33371
rect 17451 33368 17463 33371
rect 17862 33368 17868 33380
rect 17451 33340 17868 33368
rect 17451 33337 17463 33340
rect 17405 33331 17463 33337
rect 17862 33328 17868 33340
rect 17920 33328 17926 33380
rect 14645 33303 14703 33309
rect 14645 33269 14657 33303
rect 14691 33300 14703 33303
rect 14734 33300 14740 33312
rect 14691 33272 14740 33300
rect 14691 33269 14703 33272
rect 14645 33263 14703 33269
rect 14734 33260 14740 33272
rect 14792 33260 14798 33312
rect 15194 33260 15200 33312
rect 15252 33300 15258 33312
rect 16298 33300 16304 33312
rect 15252 33272 16304 33300
rect 15252 33260 15258 33272
rect 16298 33260 16304 33272
rect 16356 33260 16362 33312
rect 1104 33210 18860 33232
rect 1104 33158 3915 33210
rect 3967 33158 3979 33210
rect 4031 33158 4043 33210
rect 4095 33158 4107 33210
rect 4159 33158 4171 33210
rect 4223 33158 9846 33210
rect 9898 33158 9910 33210
rect 9962 33158 9974 33210
rect 10026 33158 10038 33210
rect 10090 33158 10102 33210
rect 10154 33158 15776 33210
rect 15828 33158 15840 33210
rect 15892 33158 15904 33210
rect 15956 33158 15968 33210
rect 16020 33158 16032 33210
rect 16084 33158 18860 33210
rect 1104 33136 18860 33158
rect 15102 33096 15108 33108
rect 15063 33068 15108 33096
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 15212 33068 16528 33096
rect 14734 32988 14740 33040
rect 14792 33028 14798 33040
rect 15212 33028 15240 33068
rect 14792 33000 15240 33028
rect 15396 33000 16436 33028
rect 14792 32988 14798 33000
rect 14550 32920 14556 32972
rect 14608 32920 14614 32972
rect 14274 32892 14280 32904
rect 14235 32864 14280 32892
rect 14274 32852 14280 32864
rect 14332 32852 14338 32904
rect 14369 32895 14427 32901
rect 14369 32861 14381 32895
rect 14415 32892 14427 32895
rect 14568 32892 14596 32920
rect 14415 32864 14596 32892
rect 14415 32861 14427 32864
rect 14369 32855 14427 32861
rect 14384 32824 14412 32855
rect 15194 32852 15200 32904
rect 15252 32892 15258 32904
rect 15396 32901 15424 33000
rect 15289 32895 15347 32901
rect 15289 32892 15301 32895
rect 15252 32864 15301 32892
rect 15252 32852 15258 32864
rect 15289 32861 15301 32864
rect 15335 32861 15347 32895
rect 15289 32855 15347 32861
rect 15381 32895 15439 32901
rect 15381 32861 15393 32895
rect 15427 32861 15439 32895
rect 15381 32855 15439 32861
rect 15473 32895 15531 32901
rect 15473 32861 15485 32895
rect 15519 32861 15531 32895
rect 15473 32855 15531 32861
rect 15565 32895 15623 32901
rect 15565 32861 15577 32895
rect 15611 32861 15623 32895
rect 16298 32892 16304 32904
rect 16259 32864 16304 32892
rect 15565 32855 15623 32861
rect 13464 32796 14412 32824
rect 14553 32827 14611 32833
rect 12710 32716 12716 32768
rect 12768 32756 12774 32768
rect 12897 32759 12955 32765
rect 12897 32756 12909 32759
rect 12768 32728 12909 32756
rect 12768 32716 12774 32728
rect 12897 32725 12909 32728
rect 12943 32725 12955 32759
rect 12897 32719 12955 32725
rect 13354 32716 13360 32768
rect 13412 32756 13418 32768
rect 13464 32765 13492 32796
rect 14553 32793 14565 32827
rect 14599 32824 14611 32827
rect 14826 32824 14832 32836
rect 14599 32796 14832 32824
rect 14599 32793 14611 32796
rect 14553 32787 14611 32793
rect 14826 32784 14832 32796
rect 14884 32824 14890 32836
rect 15488 32824 15516 32855
rect 14884 32796 15516 32824
rect 14884 32784 14890 32796
rect 13449 32759 13507 32765
rect 13449 32756 13461 32759
rect 13412 32728 13461 32756
rect 13412 32716 13418 32728
rect 13449 32725 13461 32728
rect 13495 32725 13507 32759
rect 15580 32756 15608 32855
rect 16298 32852 16304 32864
rect 16356 32852 16362 32904
rect 16408 32824 16436 33000
rect 16500 32901 16528 33068
rect 16574 33056 16580 33108
rect 16632 33096 16638 33108
rect 16850 33096 16856 33108
rect 16632 33068 16856 33096
rect 16632 33056 16638 33068
rect 16850 33056 16856 33068
rect 16908 33056 16914 33108
rect 17221 32963 17279 32969
rect 17221 32960 17233 32963
rect 16592 32932 17233 32960
rect 16485 32895 16543 32901
rect 16485 32861 16497 32895
rect 16531 32861 16543 32895
rect 16485 32855 16543 32861
rect 16592 32824 16620 32932
rect 17221 32929 17233 32932
rect 17267 32960 17279 32963
rect 17494 32960 17500 32972
rect 17267 32932 17500 32960
rect 17267 32929 17279 32932
rect 17221 32923 17279 32929
rect 17494 32920 17500 32932
rect 17552 32960 17558 32972
rect 17770 32960 17776 32972
rect 17552 32932 17776 32960
rect 17552 32920 17558 32932
rect 17770 32920 17776 32932
rect 17828 32920 17834 32972
rect 16850 32892 16856 32904
rect 16811 32864 16856 32892
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 16942 32852 16948 32904
rect 17000 32892 17006 32904
rect 17313 32895 17371 32901
rect 17313 32892 17325 32895
rect 17000 32864 17325 32892
rect 17000 32852 17006 32864
rect 17313 32861 17325 32864
rect 17359 32861 17371 32895
rect 17313 32855 17371 32861
rect 17681 32895 17739 32901
rect 17681 32861 17693 32895
rect 17727 32861 17739 32895
rect 17681 32855 17739 32861
rect 16408 32796 16620 32824
rect 17034 32756 17040 32768
rect 15580 32728 17040 32756
rect 13449 32719 13507 32725
rect 17034 32716 17040 32728
rect 17092 32716 17098 32768
rect 17310 32716 17316 32768
rect 17368 32756 17374 32768
rect 17696 32756 17724 32855
rect 17368 32728 17724 32756
rect 17368 32716 17374 32728
rect 1104 32666 18860 32688
rect 1104 32614 6880 32666
rect 6932 32614 6944 32666
rect 6996 32614 7008 32666
rect 7060 32614 7072 32666
rect 7124 32614 7136 32666
rect 7188 32614 12811 32666
rect 12863 32614 12875 32666
rect 12927 32614 12939 32666
rect 12991 32614 13003 32666
rect 13055 32614 13067 32666
rect 13119 32614 18860 32666
rect 1104 32592 18860 32614
rect 13630 32552 13636 32564
rect 13591 32524 13636 32552
rect 13630 32512 13636 32524
rect 13688 32512 13694 32564
rect 15194 32512 15200 32564
rect 15252 32552 15258 32564
rect 16117 32555 16175 32561
rect 15252 32524 16068 32552
rect 15252 32512 15258 32524
rect 15286 32484 15292 32496
rect 14292 32456 15292 32484
rect 14090 32416 14096 32428
rect 14051 32388 14096 32416
rect 14090 32376 14096 32388
rect 14148 32376 14154 32428
rect 14292 32425 14320 32456
rect 15286 32444 15292 32456
rect 15344 32444 15350 32496
rect 16040 32484 16068 32524
rect 16117 32521 16129 32555
rect 16163 32552 16175 32555
rect 16942 32552 16948 32564
rect 16163 32524 16948 32552
rect 16163 32521 16175 32524
rect 16117 32515 16175 32521
rect 16942 32512 16948 32524
rect 17000 32512 17006 32564
rect 17402 32552 17408 32564
rect 17363 32524 17408 32552
rect 17402 32512 17408 32524
rect 17460 32512 17466 32564
rect 18049 32555 18107 32561
rect 18049 32521 18061 32555
rect 18095 32552 18107 32555
rect 18138 32552 18144 32564
rect 18095 32524 18144 32552
rect 18095 32521 18107 32524
rect 18049 32515 18107 32521
rect 18138 32512 18144 32524
rect 18196 32512 18202 32564
rect 16040 32456 16712 32484
rect 14277 32419 14335 32425
rect 14277 32385 14289 32419
rect 14323 32385 14335 32419
rect 14734 32416 14740 32428
rect 14695 32388 14740 32416
rect 14277 32379 14335 32385
rect 14734 32376 14740 32388
rect 14792 32376 14798 32428
rect 14826 32376 14832 32428
rect 14884 32416 14890 32428
rect 15013 32419 15071 32425
rect 14884 32388 14977 32416
rect 14884 32376 14890 32388
rect 14936 32280 14964 32388
rect 15013 32385 15025 32419
rect 15059 32416 15071 32419
rect 15562 32416 15568 32428
rect 15059 32388 15568 32416
rect 15059 32385 15071 32388
rect 15013 32379 15071 32385
rect 15562 32376 15568 32388
rect 15620 32376 15626 32428
rect 15657 32419 15715 32425
rect 15657 32385 15669 32419
rect 15703 32416 15715 32419
rect 16574 32416 16580 32428
rect 15703 32388 16580 32416
rect 15703 32385 15715 32388
rect 15657 32379 15715 32385
rect 16574 32376 16580 32388
rect 16632 32376 16638 32428
rect 16684 32425 16712 32456
rect 17586 32444 17592 32496
rect 17644 32484 17650 32496
rect 17644 32456 18092 32484
rect 17644 32444 17650 32456
rect 16669 32419 16727 32425
rect 16669 32385 16681 32419
rect 16715 32416 16727 32419
rect 16758 32416 16764 32428
rect 16715 32388 16764 32416
rect 16715 32385 16727 32388
rect 16669 32379 16727 32385
rect 16758 32376 16764 32388
rect 16816 32376 16822 32428
rect 16850 32376 16856 32428
rect 16908 32416 16914 32428
rect 16908 32388 16953 32416
rect 16908 32376 16914 32388
rect 17034 32376 17040 32428
rect 17092 32416 17098 32428
rect 18064 32425 18092 32456
rect 17129 32419 17187 32425
rect 17129 32416 17141 32419
rect 17092 32388 17141 32416
rect 17092 32376 17098 32388
rect 17129 32385 17141 32388
rect 17175 32385 17187 32419
rect 17129 32379 17187 32385
rect 17865 32419 17923 32425
rect 17865 32385 17877 32419
rect 17911 32385 17923 32419
rect 17865 32379 17923 32385
rect 18049 32419 18107 32425
rect 18049 32385 18061 32419
rect 18095 32385 18107 32419
rect 18049 32379 18107 32385
rect 16868 32348 16896 32376
rect 15580 32320 16896 32348
rect 15580 32280 15608 32320
rect 16022 32280 16028 32292
rect 14936 32252 15608 32280
rect 15948 32252 16028 32280
rect 14093 32215 14151 32221
rect 14093 32181 14105 32215
rect 14139 32212 14151 32215
rect 15010 32212 15016 32224
rect 14139 32184 15016 32212
rect 14139 32181 14151 32184
rect 14093 32175 14151 32181
rect 15010 32172 15016 32184
rect 15068 32172 15074 32224
rect 15194 32212 15200 32224
rect 15155 32184 15200 32212
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 15948 32221 15976 32252
rect 16022 32240 16028 32252
rect 16080 32240 16086 32292
rect 16666 32240 16672 32292
rect 16724 32280 16730 32292
rect 16945 32283 17003 32289
rect 16945 32280 16957 32283
rect 16724 32252 16957 32280
rect 16724 32240 16730 32252
rect 16945 32249 16957 32252
rect 16991 32249 17003 32283
rect 16945 32243 17003 32249
rect 17037 32283 17095 32289
rect 17037 32249 17049 32283
rect 17083 32280 17095 32283
rect 17126 32280 17132 32292
rect 17083 32252 17132 32280
rect 17083 32249 17095 32252
rect 17037 32243 17095 32249
rect 17126 32240 17132 32252
rect 17184 32280 17190 32292
rect 17678 32280 17684 32292
rect 17184 32252 17684 32280
rect 17184 32240 17190 32252
rect 17678 32240 17684 32252
rect 17736 32240 17742 32292
rect 15933 32215 15991 32221
rect 15933 32181 15945 32215
rect 15979 32181 15991 32215
rect 15933 32175 15991 32181
rect 16574 32172 16580 32224
rect 16632 32212 16638 32224
rect 17880 32212 17908 32379
rect 16632 32184 17908 32212
rect 16632 32172 16638 32184
rect 1104 32122 18860 32144
rect 1104 32070 3915 32122
rect 3967 32070 3979 32122
rect 4031 32070 4043 32122
rect 4095 32070 4107 32122
rect 4159 32070 4171 32122
rect 4223 32070 9846 32122
rect 9898 32070 9910 32122
rect 9962 32070 9974 32122
rect 10026 32070 10038 32122
rect 10090 32070 10102 32122
rect 10154 32070 15776 32122
rect 15828 32070 15840 32122
rect 15892 32070 15904 32122
rect 15956 32070 15968 32122
rect 16020 32070 16032 32122
rect 16084 32070 18860 32122
rect 1104 32048 18860 32070
rect 15010 31968 15016 32020
rect 15068 32008 15074 32020
rect 15470 32008 15476 32020
rect 15068 31980 15476 32008
rect 15068 31968 15074 31980
rect 15470 31968 15476 31980
rect 15528 31968 15534 32020
rect 17034 31968 17040 32020
rect 17092 32008 17098 32020
rect 17221 32011 17279 32017
rect 17221 32008 17233 32011
rect 17092 31980 17233 32008
rect 17092 31968 17098 31980
rect 17221 31977 17233 31980
rect 17267 32008 17279 32011
rect 17494 32008 17500 32020
rect 17267 31980 17500 32008
rect 17267 31977 17279 31980
rect 17221 31971 17279 31977
rect 17494 31968 17500 31980
rect 17552 31968 17558 32020
rect 17589 31943 17647 31949
rect 17589 31940 17601 31943
rect 15396 31912 17601 31940
rect 14734 31872 14740 31884
rect 14695 31844 14740 31872
rect 14734 31832 14740 31844
rect 14792 31832 14798 31884
rect 13354 31764 13360 31816
rect 13412 31804 13418 31816
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13412 31776 14105 31804
rect 13412 31764 13418 31776
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 15396 31804 15424 31912
rect 17589 31909 17601 31912
rect 17635 31940 17647 31943
rect 17678 31940 17684 31952
rect 17635 31912 17684 31940
rect 17635 31909 17647 31912
rect 17589 31903 17647 31909
rect 17678 31900 17684 31912
rect 17736 31900 17742 31952
rect 16850 31832 16856 31884
rect 16908 31872 16914 31884
rect 16908 31844 17540 31872
rect 16908 31832 16914 31844
rect 17512 31816 17540 31844
rect 15657 31807 15715 31813
rect 15657 31804 15669 31807
rect 15396 31776 15669 31804
rect 14093 31767 14151 31773
rect 15657 31773 15669 31776
rect 15703 31773 15715 31807
rect 16393 31807 16451 31813
rect 16393 31804 16405 31807
rect 15657 31767 15715 31773
rect 16132 31776 16405 31804
rect 16132 31736 16160 31776
rect 16393 31773 16405 31776
rect 16439 31773 16451 31807
rect 16393 31767 16451 31773
rect 16758 31764 16764 31816
rect 16816 31804 16822 31816
rect 17129 31807 17187 31813
rect 17129 31804 17141 31807
rect 16816 31776 17141 31804
rect 16816 31764 16822 31776
rect 17129 31773 17141 31776
rect 17175 31804 17187 31807
rect 17310 31804 17316 31816
rect 17175 31776 17316 31804
rect 17175 31773 17187 31776
rect 17129 31767 17187 31773
rect 17310 31764 17316 31776
rect 17368 31764 17374 31816
rect 17494 31764 17500 31816
rect 17552 31764 17558 31816
rect 17402 31736 17408 31748
rect 16132 31708 17408 31736
rect 17402 31696 17408 31708
rect 17460 31696 17466 31748
rect 1104 31578 18860 31600
rect 1104 31526 6880 31578
rect 6932 31526 6944 31578
rect 6996 31526 7008 31578
rect 7060 31526 7072 31578
rect 7124 31526 7136 31578
rect 7188 31526 12811 31578
rect 12863 31526 12875 31578
rect 12927 31526 12939 31578
rect 12991 31526 13003 31578
rect 13055 31526 13067 31578
rect 13119 31526 18860 31578
rect 1104 31504 18860 31526
rect 15562 31424 15568 31476
rect 15620 31464 15626 31476
rect 16669 31467 16727 31473
rect 16669 31464 16681 31467
rect 15620 31436 16681 31464
rect 15620 31424 15626 31436
rect 16669 31433 16681 31436
rect 16715 31433 16727 31467
rect 16669 31427 16727 31433
rect 17034 31424 17040 31476
rect 17092 31424 17098 31476
rect 17954 31464 17960 31476
rect 17915 31436 17960 31464
rect 17954 31424 17960 31436
rect 18012 31424 18018 31476
rect 12710 31356 12716 31408
rect 12768 31396 12774 31408
rect 16025 31399 16083 31405
rect 16025 31396 16037 31399
rect 12768 31368 16037 31396
rect 12768 31356 12774 31368
rect 16025 31365 16037 31368
rect 16071 31396 16083 31399
rect 16574 31396 16580 31408
rect 16071 31368 16580 31396
rect 16071 31365 16083 31368
rect 16025 31359 16083 31365
rect 16574 31356 16580 31368
rect 16632 31356 16638 31408
rect 17052 31396 17080 31424
rect 17052 31368 17632 31396
rect 14090 31288 14096 31340
rect 14148 31328 14154 31340
rect 15381 31331 15439 31337
rect 15381 31328 15393 31331
rect 14148 31300 15393 31328
rect 14148 31288 14154 31300
rect 15381 31297 15393 31300
rect 15427 31297 15439 31331
rect 15381 31291 15439 31297
rect 16482 31288 16488 31340
rect 16540 31328 16546 31340
rect 16853 31331 16911 31337
rect 16853 31328 16865 31331
rect 16540 31300 16865 31328
rect 16540 31288 16546 31300
rect 16853 31297 16865 31300
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 16942 31288 16948 31340
rect 17000 31328 17006 31340
rect 17037 31331 17095 31337
rect 17037 31328 17049 31331
rect 17000 31300 17049 31328
rect 17000 31288 17006 31300
rect 17037 31297 17049 31300
rect 17083 31297 17095 31331
rect 17037 31291 17095 31297
rect 17126 31288 17132 31340
rect 17184 31328 17190 31340
rect 17604 31337 17632 31368
rect 17589 31331 17647 31337
rect 17184 31300 17229 31328
rect 17184 31288 17190 31300
rect 17589 31297 17601 31331
rect 17635 31297 17647 31331
rect 17589 31291 17647 31297
rect 17678 31288 17684 31340
rect 17736 31328 17742 31340
rect 17736 31300 17781 31328
rect 17736 31288 17742 31300
rect 15197 31263 15255 31269
rect 15197 31229 15209 31263
rect 15243 31260 15255 31263
rect 15286 31260 15292 31272
rect 15243 31232 15292 31260
rect 15243 31229 15255 31232
rect 15197 31223 15255 31229
rect 15286 31220 15292 31232
rect 15344 31220 15350 31272
rect 15565 31195 15623 31201
rect 15565 31161 15577 31195
rect 15611 31192 15623 31195
rect 16114 31192 16120 31204
rect 15611 31164 16120 31192
rect 15611 31161 15623 31164
rect 15565 31155 15623 31161
rect 16114 31152 16120 31164
rect 16172 31152 16178 31204
rect 16666 31084 16672 31136
rect 16724 31124 16730 31136
rect 17589 31127 17647 31133
rect 17589 31124 17601 31127
rect 16724 31096 17601 31124
rect 16724 31084 16730 31096
rect 17589 31093 17601 31096
rect 17635 31093 17647 31127
rect 17589 31087 17647 31093
rect 1104 31034 18860 31056
rect 1104 30982 3915 31034
rect 3967 30982 3979 31034
rect 4031 30982 4043 31034
rect 4095 30982 4107 31034
rect 4159 30982 4171 31034
rect 4223 30982 9846 31034
rect 9898 30982 9910 31034
rect 9962 30982 9974 31034
rect 10026 30982 10038 31034
rect 10090 30982 10102 31034
rect 10154 30982 15776 31034
rect 15828 30982 15840 31034
rect 15892 30982 15904 31034
rect 15956 30982 15968 31034
rect 16020 30982 16032 31034
rect 16084 30982 18860 31034
rect 1104 30960 18860 30982
rect 17402 30920 17408 30932
rect 17363 30892 17408 30920
rect 17402 30880 17408 30892
rect 17460 30880 17466 30932
rect 15194 30812 15200 30864
rect 15252 30852 15258 30864
rect 16853 30855 16911 30861
rect 15252 30824 16712 30852
rect 15252 30812 15258 30824
rect 1394 30716 1400 30728
rect 1355 30688 1400 30716
rect 1394 30676 1400 30688
rect 1452 30676 1458 30728
rect 1673 30719 1731 30725
rect 1673 30685 1685 30719
rect 1719 30716 1731 30719
rect 14090 30716 14096 30728
rect 1719 30688 14096 30716
rect 1719 30685 1731 30688
rect 1673 30679 1731 30685
rect 14090 30676 14096 30688
rect 14148 30676 14154 30728
rect 15470 30676 15476 30728
rect 15528 30716 15534 30728
rect 15841 30719 15899 30725
rect 15841 30716 15853 30719
rect 15528 30688 15853 30716
rect 15528 30676 15534 30688
rect 15841 30685 15853 30688
rect 15887 30685 15899 30719
rect 16022 30716 16028 30728
rect 15983 30688 16028 30716
rect 15841 30679 15899 30685
rect 16022 30676 16028 30688
rect 16080 30676 16086 30728
rect 16684 30725 16712 30824
rect 16853 30821 16865 30855
rect 16899 30852 16911 30855
rect 18138 30852 18144 30864
rect 16899 30824 18144 30852
rect 16899 30821 16911 30824
rect 16853 30815 16911 30821
rect 18138 30812 18144 30824
rect 18196 30812 18202 30864
rect 17770 30784 17776 30796
rect 17328 30756 17776 30784
rect 17328 30725 17356 30756
rect 17770 30744 17776 30756
rect 17828 30744 17834 30796
rect 16577 30719 16635 30725
rect 16577 30716 16589 30719
rect 16500 30688 16589 30716
rect 16500 30648 16528 30688
rect 16577 30685 16589 30688
rect 16623 30685 16635 30719
rect 16577 30679 16635 30685
rect 16669 30719 16727 30725
rect 16669 30685 16681 30719
rect 16715 30685 16727 30719
rect 16669 30679 16727 30685
rect 17313 30719 17371 30725
rect 17313 30685 17325 30719
rect 17359 30685 17371 30719
rect 17494 30716 17500 30728
rect 17455 30688 17500 30716
rect 17313 30679 17371 30685
rect 17328 30648 17356 30679
rect 17494 30676 17500 30688
rect 17552 30676 17558 30728
rect 16500 30620 17356 30648
rect 15746 30540 15752 30592
rect 15804 30580 15810 30592
rect 15933 30583 15991 30589
rect 15933 30580 15945 30583
rect 15804 30552 15945 30580
rect 15804 30540 15810 30552
rect 15933 30549 15945 30552
rect 15979 30549 15991 30583
rect 15933 30543 15991 30549
rect 1104 30490 18860 30512
rect 1104 30438 6880 30490
rect 6932 30438 6944 30490
rect 6996 30438 7008 30490
rect 7060 30438 7072 30490
rect 7124 30438 7136 30490
rect 7188 30438 12811 30490
rect 12863 30438 12875 30490
rect 12927 30438 12939 30490
rect 12991 30438 13003 30490
rect 13055 30438 13067 30490
rect 13119 30438 18860 30490
rect 1104 30416 18860 30438
rect 1394 30376 1400 30388
rect 1355 30348 1400 30376
rect 1394 30336 1400 30348
rect 1452 30336 1458 30388
rect 17310 30376 17316 30388
rect 17271 30348 17316 30376
rect 17310 30336 17316 30348
rect 17368 30336 17374 30388
rect 15378 30268 15384 30320
rect 15436 30308 15442 30320
rect 16761 30311 16819 30317
rect 16761 30308 16773 30311
rect 15436 30280 16773 30308
rect 15436 30268 15442 30280
rect 16761 30277 16773 30280
rect 16807 30277 16819 30311
rect 16761 30271 16819 30277
rect 17328 30280 18092 30308
rect 15746 30240 15752 30252
rect 15707 30212 15752 30240
rect 15746 30200 15752 30212
rect 15804 30200 15810 30252
rect 15841 30243 15899 30249
rect 15841 30209 15853 30243
rect 15887 30209 15899 30243
rect 15841 30203 15899 30209
rect 15102 30132 15108 30184
rect 15160 30172 15166 30184
rect 15856 30172 15884 30203
rect 16022 30200 16028 30252
rect 16080 30240 16086 30252
rect 16669 30243 16727 30249
rect 16669 30240 16681 30243
rect 16080 30212 16681 30240
rect 16080 30200 16086 30212
rect 16669 30209 16681 30212
rect 16715 30209 16727 30243
rect 16669 30203 16727 30209
rect 16853 30243 16911 30249
rect 16853 30209 16865 30243
rect 16899 30240 16911 30243
rect 17126 30240 17132 30252
rect 16899 30212 17132 30240
rect 16899 30209 16911 30212
rect 16853 30203 16911 30209
rect 15160 30144 15884 30172
rect 15160 30132 15166 30144
rect 16025 30107 16083 30113
rect 16025 30073 16037 30107
rect 16071 30104 16083 30107
rect 16868 30104 16896 30203
rect 17126 30200 17132 30212
rect 17184 30200 17190 30252
rect 17328 30249 17356 30280
rect 18064 30252 18092 30280
rect 17313 30243 17371 30249
rect 17313 30209 17325 30243
rect 17359 30209 17371 30243
rect 17313 30203 17371 30209
rect 17497 30243 17555 30249
rect 17497 30209 17509 30243
rect 17543 30240 17555 30243
rect 17862 30240 17868 30252
rect 17543 30212 17868 30240
rect 17543 30209 17555 30212
rect 17497 30203 17555 30209
rect 17862 30200 17868 30212
rect 17920 30240 17926 30252
rect 17957 30243 18015 30249
rect 17957 30240 17969 30243
rect 17920 30212 17969 30240
rect 17920 30200 17926 30212
rect 17957 30209 17969 30212
rect 18003 30209 18015 30243
rect 17957 30203 18015 30209
rect 18046 30200 18052 30252
rect 18104 30240 18110 30252
rect 18141 30243 18199 30249
rect 18141 30240 18153 30243
rect 18104 30212 18153 30240
rect 18104 30200 18110 30212
rect 18141 30209 18153 30212
rect 18187 30209 18199 30243
rect 18141 30203 18199 30209
rect 16071 30076 16896 30104
rect 16071 30073 16083 30076
rect 16025 30067 16083 30073
rect 17586 30064 17592 30116
rect 17644 30104 17650 30116
rect 17957 30107 18015 30113
rect 17957 30104 17969 30107
rect 17644 30076 17969 30104
rect 17644 30064 17650 30076
rect 17957 30073 17969 30076
rect 18003 30073 18015 30107
rect 17957 30067 18015 30073
rect 1104 29946 18860 29968
rect 1104 29894 3915 29946
rect 3967 29894 3979 29946
rect 4031 29894 4043 29946
rect 4095 29894 4107 29946
rect 4159 29894 4171 29946
rect 4223 29894 9846 29946
rect 9898 29894 9910 29946
rect 9962 29894 9974 29946
rect 10026 29894 10038 29946
rect 10090 29894 10102 29946
rect 10154 29894 15776 29946
rect 15828 29894 15840 29946
rect 15892 29894 15904 29946
rect 15956 29894 15968 29946
rect 16020 29894 16032 29946
rect 16084 29894 18860 29946
rect 1104 29872 18860 29894
rect 14366 29656 14372 29708
rect 14424 29696 14430 29708
rect 15102 29696 15108 29708
rect 14424 29668 15108 29696
rect 14424 29656 14430 29668
rect 15102 29656 15108 29668
rect 15160 29696 15166 29708
rect 15160 29668 16068 29696
rect 15160 29656 15166 29668
rect 15654 29588 15660 29640
rect 15712 29628 15718 29640
rect 16040 29637 16068 29668
rect 15841 29631 15899 29637
rect 15841 29628 15853 29631
rect 15712 29600 15853 29628
rect 15712 29588 15718 29600
rect 15841 29597 15853 29600
rect 15887 29597 15899 29631
rect 15841 29591 15899 29597
rect 16025 29631 16083 29637
rect 16025 29597 16037 29631
rect 16071 29597 16083 29631
rect 16025 29591 16083 29597
rect 17126 29588 17132 29640
rect 17184 29628 17190 29640
rect 17773 29631 17831 29637
rect 17773 29628 17785 29631
rect 17184 29600 17785 29628
rect 17184 29588 17190 29600
rect 17773 29597 17785 29600
rect 17819 29597 17831 29631
rect 17773 29591 17831 29597
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29597 18015 29631
rect 17957 29591 18015 29597
rect 15933 29563 15991 29569
rect 15933 29529 15945 29563
rect 15979 29560 15991 29563
rect 17972 29560 18000 29591
rect 15979 29532 18000 29560
rect 15979 29529 15991 29532
rect 15933 29523 15991 29529
rect 13630 29452 13636 29504
rect 13688 29492 13694 29504
rect 15562 29492 15568 29504
rect 13688 29464 15568 29492
rect 13688 29452 13694 29464
rect 15562 29452 15568 29464
rect 15620 29452 15626 29504
rect 17954 29452 17960 29504
rect 18012 29492 18018 29504
rect 18049 29495 18107 29501
rect 18049 29492 18061 29495
rect 18012 29464 18061 29492
rect 18012 29452 18018 29464
rect 18049 29461 18061 29464
rect 18095 29461 18107 29495
rect 18049 29455 18107 29461
rect 1104 29402 18860 29424
rect 1104 29350 6880 29402
rect 6932 29350 6944 29402
rect 6996 29350 7008 29402
rect 7060 29350 7072 29402
rect 7124 29350 7136 29402
rect 7188 29350 12811 29402
rect 12863 29350 12875 29402
rect 12927 29350 12939 29402
rect 12991 29350 13003 29402
rect 13055 29350 13067 29402
rect 13119 29350 18860 29402
rect 1104 29328 18860 29350
rect 1104 28858 18860 28880
rect 1104 28806 3915 28858
rect 3967 28806 3979 28858
rect 4031 28806 4043 28858
rect 4095 28806 4107 28858
rect 4159 28806 4171 28858
rect 4223 28806 9846 28858
rect 9898 28806 9910 28858
rect 9962 28806 9974 28858
rect 10026 28806 10038 28858
rect 10090 28806 10102 28858
rect 10154 28806 15776 28858
rect 15828 28806 15840 28858
rect 15892 28806 15904 28858
rect 15956 28806 15968 28858
rect 16020 28806 16032 28858
rect 16084 28806 18860 28858
rect 1104 28784 18860 28806
rect 16206 28704 16212 28756
rect 16264 28744 16270 28756
rect 17957 28747 18015 28753
rect 17957 28744 17969 28747
rect 16264 28716 17969 28744
rect 16264 28704 16270 28716
rect 17957 28713 17969 28716
rect 18003 28713 18015 28747
rect 17957 28707 18015 28713
rect 17497 28543 17555 28549
rect 17497 28509 17509 28543
rect 17543 28540 17555 28543
rect 18138 28540 18144 28552
rect 17543 28512 18144 28540
rect 17543 28509 17555 28512
rect 17497 28503 17555 28509
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 1104 28314 18860 28336
rect 1104 28262 6880 28314
rect 6932 28262 6944 28314
rect 6996 28262 7008 28314
rect 7060 28262 7072 28314
rect 7124 28262 7136 28314
rect 7188 28262 12811 28314
rect 12863 28262 12875 28314
rect 12927 28262 12939 28314
rect 12991 28262 13003 28314
rect 13055 28262 13067 28314
rect 13119 28262 18860 28314
rect 1104 28240 18860 28262
rect 1104 27770 18860 27792
rect 1104 27718 3915 27770
rect 3967 27718 3979 27770
rect 4031 27718 4043 27770
rect 4095 27718 4107 27770
rect 4159 27718 4171 27770
rect 4223 27718 9846 27770
rect 9898 27718 9910 27770
rect 9962 27718 9974 27770
rect 10026 27718 10038 27770
rect 10090 27718 10102 27770
rect 10154 27718 15776 27770
rect 15828 27718 15840 27770
rect 15892 27718 15904 27770
rect 15956 27718 15968 27770
rect 16020 27718 16032 27770
rect 16084 27718 18860 27770
rect 1104 27696 18860 27718
rect 1104 27226 18860 27248
rect 1104 27174 6880 27226
rect 6932 27174 6944 27226
rect 6996 27174 7008 27226
rect 7060 27174 7072 27226
rect 7124 27174 7136 27226
rect 7188 27174 12811 27226
rect 12863 27174 12875 27226
rect 12927 27174 12939 27226
rect 12991 27174 13003 27226
rect 13055 27174 13067 27226
rect 13119 27174 18860 27226
rect 1104 27152 18860 27174
rect 1104 26682 18860 26704
rect 1104 26630 3915 26682
rect 3967 26630 3979 26682
rect 4031 26630 4043 26682
rect 4095 26630 4107 26682
rect 4159 26630 4171 26682
rect 4223 26630 9846 26682
rect 9898 26630 9910 26682
rect 9962 26630 9974 26682
rect 10026 26630 10038 26682
rect 10090 26630 10102 26682
rect 10154 26630 15776 26682
rect 15828 26630 15840 26682
rect 15892 26630 15904 26682
rect 15956 26630 15968 26682
rect 16020 26630 16032 26682
rect 16084 26630 18860 26682
rect 1104 26608 18860 26630
rect 1104 26138 18860 26160
rect 1104 26086 6880 26138
rect 6932 26086 6944 26138
rect 6996 26086 7008 26138
rect 7060 26086 7072 26138
rect 7124 26086 7136 26138
rect 7188 26086 12811 26138
rect 12863 26086 12875 26138
rect 12927 26086 12939 26138
rect 12991 26086 13003 26138
rect 13055 26086 13067 26138
rect 13119 26086 18860 26138
rect 1104 26064 18860 26086
rect 14366 26024 14372 26036
rect 14327 25996 14372 26024
rect 14366 25984 14372 25996
rect 14424 25984 14430 26036
rect 13630 25848 13636 25900
rect 13688 25888 13694 25900
rect 14093 25891 14151 25897
rect 14093 25888 14105 25891
rect 13688 25860 14105 25888
rect 13688 25848 13694 25860
rect 14093 25857 14105 25860
rect 14139 25857 14151 25891
rect 14093 25851 14151 25857
rect 13446 25780 13452 25832
rect 13504 25820 13510 25832
rect 13725 25823 13783 25829
rect 13725 25820 13737 25823
rect 13504 25792 13737 25820
rect 13504 25780 13510 25792
rect 13725 25789 13737 25792
rect 13771 25789 13783 25823
rect 13725 25783 13783 25789
rect 14182 25780 14188 25832
rect 14240 25820 14246 25832
rect 14240 25792 14285 25820
rect 14240 25780 14246 25792
rect 1104 25594 18860 25616
rect 1104 25542 3915 25594
rect 3967 25542 3979 25594
rect 4031 25542 4043 25594
rect 4095 25542 4107 25594
rect 4159 25542 4171 25594
rect 4223 25542 9846 25594
rect 9898 25542 9910 25594
rect 9962 25542 9974 25594
rect 10026 25542 10038 25594
rect 10090 25542 10102 25594
rect 10154 25542 15776 25594
rect 15828 25542 15840 25594
rect 15892 25542 15904 25594
rect 15956 25542 15968 25594
rect 16020 25542 16032 25594
rect 16084 25542 18860 25594
rect 1104 25520 18860 25542
rect 13170 25480 13176 25492
rect 13131 25452 13176 25480
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25276 1731 25279
rect 11146 25276 11152 25288
rect 1719 25248 11152 25276
rect 1719 25245 1731 25248
rect 1673 25239 1731 25245
rect 11146 25236 11152 25248
rect 11204 25236 11210 25288
rect 1486 25140 1492 25152
rect 1447 25112 1492 25140
rect 1486 25100 1492 25112
rect 1544 25100 1550 25152
rect 1104 25050 18860 25072
rect 1104 24998 6880 25050
rect 6932 24998 6944 25050
rect 6996 24998 7008 25050
rect 7060 24998 7072 25050
rect 7124 24998 7136 25050
rect 7188 24998 12811 25050
rect 12863 24998 12875 25050
rect 12927 24998 12939 25050
rect 12991 24998 13003 25050
rect 13055 24998 13067 25050
rect 13119 24998 18860 25050
rect 1104 24976 18860 24998
rect 12805 24871 12863 24877
rect 12805 24837 12817 24871
rect 12851 24868 12863 24871
rect 13170 24868 13176 24880
rect 12851 24840 13176 24868
rect 12851 24837 12863 24840
rect 12805 24831 12863 24837
rect 13170 24828 13176 24840
rect 13228 24828 13234 24880
rect 1670 24760 1676 24812
rect 1728 24800 1734 24812
rect 12526 24800 12532 24812
rect 1728 24772 12532 24800
rect 1728 24760 1734 24772
rect 12526 24760 12532 24772
rect 12584 24800 12590 24812
rect 12621 24803 12679 24809
rect 12621 24800 12633 24803
rect 12584 24772 12633 24800
rect 12584 24760 12590 24772
rect 12621 24769 12633 24772
rect 12667 24769 12679 24803
rect 13446 24800 13452 24812
rect 13407 24772 13452 24800
rect 12621 24763 12679 24769
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 14182 24800 14188 24812
rect 13679 24772 14188 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 12989 24735 13047 24741
rect 12989 24701 13001 24735
rect 13035 24732 13047 24735
rect 13648 24732 13676 24763
rect 14182 24760 14188 24772
rect 14240 24760 14246 24812
rect 13035 24704 13676 24732
rect 13035 24701 13047 24704
rect 12989 24695 13047 24701
rect 13538 24596 13544 24608
rect 13499 24568 13544 24596
rect 13538 24556 13544 24568
rect 13596 24556 13602 24608
rect 1104 24506 18860 24528
rect 1104 24454 3915 24506
rect 3967 24454 3979 24506
rect 4031 24454 4043 24506
rect 4095 24454 4107 24506
rect 4159 24454 4171 24506
rect 4223 24454 9846 24506
rect 9898 24454 9910 24506
rect 9962 24454 9974 24506
rect 10026 24454 10038 24506
rect 10090 24454 10102 24506
rect 10154 24454 15776 24506
rect 15828 24454 15840 24506
rect 15892 24454 15904 24506
rect 15956 24454 15968 24506
rect 16020 24454 16032 24506
rect 16084 24454 18860 24506
rect 1104 24432 18860 24454
rect 12621 24395 12679 24401
rect 12621 24361 12633 24395
rect 12667 24392 12679 24395
rect 13446 24392 13452 24404
rect 12667 24364 13452 24392
rect 12667 24361 12679 24364
rect 12621 24355 12679 24361
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 11146 24324 11152 24336
rect 11107 24296 11152 24324
rect 11146 24284 11152 24296
rect 11204 24284 11210 24336
rect 13170 24324 13176 24336
rect 13131 24296 13176 24324
rect 13170 24284 13176 24296
rect 13228 24284 13234 24336
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 13538 24256 13544 24268
rect 11655 24228 13544 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 13538 24216 13544 24228
rect 13596 24216 13602 24268
rect 11517 24191 11575 24197
rect 11517 24157 11529 24191
rect 11563 24157 11575 24191
rect 12526 24188 12532 24200
rect 12487 24160 12532 24188
rect 11517 24151 11575 24157
rect 11532 24120 11560 24151
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 12713 24191 12771 24197
rect 12713 24157 12725 24191
rect 12759 24188 12771 24191
rect 13170 24188 13176 24200
rect 12759 24160 13176 24188
rect 12759 24157 12771 24160
rect 12713 24151 12771 24157
rect 13170 24148 13176 24160
rect 13228 24148 13234 24200
rect 13630 24120 13636 24132
rect 11532 24092 13636 24120
rect 13630 24080 13636 24092
rect 13688 24080 13694 24132
rect 1104 23962 18860 23984
rect 1104 23910 6880 23962
rect 6932 23910 6944 23962
rect 6996 23910 7008 23962
rect 7060 23910 7072 23962
rect 7124 23910 7136 23962
rect 7188 23910 12811 23962
rect 12863 23910 12875 23962
rect 12927 23910 12939 23962
rect 12991 23910 13003 23962
rect 13055 23910 13067 23962
rect 13119 23910 18860 23962
rect 1104 23888 18860 23910
rect 1104 23418 18860 23440
rect 1104 23366 3915 23418
rect 3967 23366 3979 23418
rect 4031 23366 4043 23418
rect 4095 23366 4107 23418
rect 4159 23366 4171 23418
rect 4223 23366 9846 23418
rect 9898 23366 9910 23418
rect 9962 23366 9974 23418
rect 10026 23366 10038 23418
rect 10090 23366 10102 23418
rect 10154 23366 15776 23418
rect 15828 23366 15840 23418
rect 15892 23366 15904 23418
rect 15956 23366 15968 23418
rect 16020 23366 16032 23418
rect 16084 23366 18860 23418
rect 1104 23344 18860 23366
rect 1104 22874 18860 22896
rect 1104 22822 6880 22874
rect 6932 22822 6944 22874
rect 6996 22822 7008 22874
rect 7060 22822 7072 22874
rect 7124 22822 7136 22874
rect 7188 22822 12811 22874
rect 12863 22822 12875 22874
rect 12927 22822 12939 22874
rect 12991 22822 13003 22874
rect 13055 22822 13067 22874
rect 13119 22822 18860 22874
rect 1104 22800 18860 22822
rect 1104 22330 18860 22352
rect 1104 22278 3915 22330
rect 3967 22278 3979 22330
rect 4031 22278 4043 22330
rect 4095 22278 4107 22330
rect 4159 22278 4171 22330
rect 4223 22278 9846 22330
rect 9898 22278 9910 22330
rect 9962 22278 9974 22330
rect 10026 22278 10038 22330
rect 10090 22278 10102 22330
rect 10154 22278 15776 22330
rect 15828 22278 15840 22330
rect 15892 22278 15904 22330
rect 15956 22278 15968 22330
rect 16020 22278 16032 22330
rect 16084 22278 18860 22330
rect 1104 22256 18860 22278
rect 13541 22083 13599 22089
rect 13541 22049 13553 22083
rect 13587 22080 13599 22083
rect 13630 22080 13636 22092
rect 13587 22052 13636 22080
rect 13587 22049 13599 22052
rect 13541 22043 13599 22049
rect 13630 22040 13636 22052
rect 13688 22040 13694 22092
rect 13998 22040 14004 22092
rect 14056 22080 14062 22092
rect 14093 22083 14151 22089
rect 14093 22080 14105 22083
rect 14056 22052 14105 22080
rect 14056 22040 14062 22052
rect 14093 22049 14105 22052
rect 14139 22049 14151 22083
rect 14093 22043 14151 22049
rect 13265 22015 13323 22021
rect 13265 21981 13277 22015
rect 13311 21981 13323 22015
rect 13265 21975 13323 21981
rect 13357 22015 13415 22021
rect 13357 21981 13369 22015
rect 13403 22012 13415 22015
rect 13446 22012 13452 22024
rect 13403 21984 13452 22012
rect 13403 21981 13415 21984
rect 13357 21975 13415 21981
rect 13280 21944 13308 21975
rect 13446 21972 13452 21984
rect 13504 21972 13510 22024
rect 14016 21944 14044 22040
rect 17497 22015 17555 22021
rect 17497 21981 17509 22015
rect 17543 22012 17555 22015
rect 18138 22012 18144 22024
rect 17543 21984 18144 22012
rect 17543 21981 17555 21984
rect 17497 21975 17555 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 13280 21916 14044 21944
rect 12897 21879 12955 21885
rect 12897 21845 12909 21879
rect 12943 21876 12955 21879
rect 13262 21876 13268 21888
rect 12943 21848 13268 21876
rect 12943 21845 12955 21848
rect 12897 21839 12955 21845
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 17957 21879 18015 21885
rect 17957 21845 17969 21879
rect 18003 21876 18015 21879
rect 18046 21876 18052 21888
rect 18003 21848 18052 21876
rect 18003 21845 18015 21848
rect 17957 21839 18015 21845
rect 18046 21836 18052 21848
rect 18104 21836 18110 21888
rect 1104 21786 18860 21808
rect 1104 21734 6880 21786
rect 6932 21734 6944 21786
rect 6996 21734 7008 21786
rect 7060 21734 7072 21786
rect 7124 21734 7136 21786
rect 7188 21734 12811 21786
rect 12863 21734 12875 21786
rect 12927 21734 12939 21786
rect 12991 21734 13003 21786
rect 13055 21734 13067 21786
rect 13119 21734 18860 21786
rect 1104 21712 18860 21734
rect 1104 21242 18860 21264
rect 1104 21190 3915 21242
rect 3967 21190 3979 21242
rect 4031 21190 4043 21242
rect 4095 21190 4107 21242
rect 4159 21190 4171 21242
rect 4223 21190 9846 21242
rect 9898 21190 9910 21242
rect 9962 21190 9974 21242
rect 10026 21190 10038 21242
rect 10090 21190 10102 21242
rect 10154 21190 15776 21242
rect 15828 21190 15840 21242
rect 15892 21190 15904 21242
rect 15956 21190 15968 21242
rect 16020 21190 16032 21242
rect 16084 21190 18860 21242
rect 1104 21168 18860 21190
rect 1104 20698 18860 20720
rect 1104 20646 6880 20698
rect 6932 20646 6944 20698
rect 6996 20646 7008 20698
rect 7060 20646 7072 20698
rect 7124 20646 7136 20698
rect 7188 20646 12811 20698
rect 12863 20646 12875 20698
rect 12927 20646 12939 20698
rect 12991 20646 13003 20698
rect 13055 20646 13067 20698
rect 13119 20646 18860 20698
rect 1104 20624 18860 20646
rect 13262 20448 13268 20460
rect 13223 20420 13268 20448
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13446 20448 13452 20460
rect 13407 20420 13452 20448
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13357 20247 13415 20253
rect 13357 20213 13369 20247
rect 13403 20244 13415 20247
rect 15010 20244 15016 20256
rect 13403 20216 15016 20244
rect 13403 20213 13415 20216
rect 13357 20207 13415 20213
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 1104 20154 18860 20176
rect 1104 20102 3915 20154
rect 3967 20102 3979 20154
rect 4031 20102 4043 20154
rect 4095 20102 4107 20154
rect 4159 20102 4171 20154
rect 4223 20102 9846 20154
rect 9898 20102 9910 20154
rect 9962 20102 9974 20154
rect 10026 20102 10038 20154
rect 10090 20102 10102 20154
rect 10154 20102 15776 20154
rect 15828 20102 15840 20154
rect 15892 20102 15904 20154
rect 15956 20102 15968 20154
rect 16020 20102 16032 20154
rect 16084 20102 18860 20154
rect 1104 20080 18860 20102
rect 1670 19904 1676 19916
rect 1631 19876 1676 19904
rect 1670 19864 1676 19876
rect 1728 19864 1734 19916
rect 1394 19836 1400 19848
rect 1355 19808 1400 19836
rect 1394 19796 1400 19808
rect 1452 19796 1458 19848
rect 1104 19610 18860 19632
rect 1104 19558 6880 19610
rect 6932 19558 6944 19610
rect 6996 19558 7008 19610
rect 7060 19558 7072 19610
rect 7124 19558 7136 19610
rect 7188 19558 12811 19610
rect 12863 19558 12875 19610
rect 12927 19558 12939 19610
rect 12991 19558 13003 19610
rect 13055 19558 13067 19610
rect 13119 19558 18860 19610
rect 1104 19536 18860 19558
rect 1394 19428 1400 19440
rect 1355 19400 1400 19428
rect 1394 19388 1400 19400
rect 1452 19388 1458 19440
rect 15289 19363 15347 19369
rect 15289 19360 15301 19363
rect 14936 19332 15301 19360
rect 13998 19252 14004 19304
rect 14056 19292 14062 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 14056 19264 14473 19292
rect 14056 19252 14062 19264
rect 14461 19261 14473 19264
rect 14507 19292 14519 19295
rect 14936 19292 14964 19332
rect 15289 19329 15301 19332
rect 15335 19329 15347 19363
rect 15289 19323 15347 19329
rect 14507 19264 14964 19292
rect 14507 19261 14519 19264
rect 14461 19255 14519 19261
rect 15010 19252 15016 19304
rect 15068 19292 15074 19304
rect 15197 19295 15255 19301
rect 15197 19292 15209 19295
rect 15068 19264 15209 19292
rect 15068 19252 15074 19264
rect 15197 19261 15209 19264
rect 15243 19261 15255 19295
rect 16114 19292 16120 19304
rect 16075 19264 16120 19292
rect 15197 19255 15255 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 1104 19066 18860 19088
rect 1104 19014 3915 19066
rect 3967 19014 3979 19066
rect 4031 19014 4043 19066
rect 4095 19014 4107 19066
rect 4159 19014 4171 19066
rect 4223 19014 9846 19066
rect 9898 19014 9910 19066
rect 9962 19014 9974 19066
rect 10026 19014 10038 19066
rect 10090 19014 10102 19066
rect 10154 19014 15776 19066
rect 15828 19014 15840 19066
rect 15892 19014 15904 19066
rect 15956 19014 15968 19066
rect 16020 19014 16032 19066
rect 16084 19014 18860 19066
rect 1104 18992 18860 19014
rect 1104 18522 18860 18544
rect 1104 18470 6880 18522
rect 6932 18470 6944 18522
rect 6996 18470 7008 18522
rect 7060 18470 7072 18522
rect 7124 18470 7136 18522
rect 7188 18470 12811 18522
rect 12863 18470 12875 18522
rect 12927 18470 12939 18522
rect 12991 18470 13003 18522
rect 13055 18470 13067 18522
rect 13119 18470 18860 18522
rect 1104 18448 18860 18470
rect 10965 18411 11023 18417
rect 10965 18377 10977 18411
rect 11011 18408 11023 18411
rect 11885 18411 11943 18417
rect 11011 18380 11836 18408
rect 11011 18377 11023 18380
rect 10965 18371 11023 18377
rect 11808 18340 11836 18380
rect 11885 18377 11897 18411
rect 11931 18408 11943 18411
rect 13446 18408 13452 18420
rect 11931 18380 13452 18408
rect 11931 18377 11943 18380
rect 11885 18371 11943 18377
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 13262 18340 13268 18352
rect 10796 18312 11376 18340
rect 11808 18312 13268 18340
rect 10796 18281 10824 18312
rect 11348 18284 11376 18312
rect 13262 18300 13268 18312
rect 13320 18300 13326 18352
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10367 18244 10793 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 10965 18275 11023 18281
rect 10965 18241 10977 18275
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 10980 18204 11008 18235
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11388 18244 11529 18272
rect 11388 18232 11394 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18241 11759 18275
rect 11701 18235 11759 18241
rect 11716 18204 11744 18235
rect 8352 18176 11744 18204
rect 8352 18164 8358 18176
rect 1104 17978 18860 18000
rect 1104 17926 3915 17978
rect 3967 17926 3979 17978
rect 4031 17926 4043 17978
rect 4095 17926 4107 17978
rect 4159 17926 4171 17978
rect 4223 17926 9846 17978
rect 9898 17926 9910 17978
rect 9962 17926 9974 17978
rect 10026 17926 10038 17978
rect 10090 17926 10102 17978
rect 10154 17926 15776 17978
rect 15828 17926 15840 17978
rect 15892 17926 15904 17978
rect 15956 17926 15968 17978
rect 16020 17926 16032 17978
rect 16084 17926 18860 17978
rect 1104 17904 18860 17926
rect 11330 17524 11336 17536
rect 11291 17496 11336 17524
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 1104 17434 18860 17456
rect 1104 17382 6880 17434
rect 6932 17382 6944 17434
rect 6996 17382 7008 17434
rect 7060 17382 7072 17434
rect 7124 17382 7136 17434
rect 7188 17382 12811 17434
rect 12863 17382 12875 17434
rect 12927 17382 12939 17434
rect 12991 17382 13003 17434
rect 13055 17382 13067 17434
rect 13119 17382 18860 17434
rect 1104 17360 18860 17382
rect 1104 16890 18860 16912
rect 1104 16838 3915 16890
rect 3967 16838 3979 16890
rect 4031 16838 4043 16890
rect 4095 16838 4107 16890
rect 4159 16838 4171 16890
rect 4223 16838 9846 16890
rect 9898 16838 9910 16890
rect 9962 16838 9974 16890
rect 10026 16838 10038 16890
rect 10090 16838 10102 16890
rect 10154 16838 15776 16890
rect 15828 16838 15840 16890
rect 15892 16838 15904 16890
rect 15956 16838 15968 16890
rect 16020 16838 16032 16890
rect 16084 16838 18860 16890
rect 1104 16816 18860 16838
rect 1104 16346 18860 16368
rect 1104 16294 6880 16346
rect 6932 16294 6944 16346
rect 6996 16294 7008 16346
rect 7060 16294 7072 16346
rect 7124 16294 7136 16346
rect 7188 16294 12811 16346
rect 12863 16294 12875 16346
rect 12927 16294 12939 16346
rect 12991 16294 13003 16346
rect 13055 16294 13067 16346
rect 13119 16294 18860 16346
rect 1104 16272 18860 16294
rect 17862 16096 17868 16108
rect 17823 16068 17868 16096
rect 17862 16056 17868 16068
rect 17920 16056 17926 16108
rect 18138 16028 18144 16040
rect 18099 16000 18144 16028
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 1104 15802 18860 15824
rect 1104 15750 3915 15802
rect 3967 15750 3979 15802
rect 4031 15750 4043 15802
rect 4095 15750 4107 15802
rect 4159 15750 4171 15802
rect 4223 15750 9846 15802
rect 9898 15750 9910 15802
rect 9962 15750 9974 15802
rect 10026 15750 10038 15802
rect 10090 15750 10102 15802
rect 10154 15750 15776 15802
rect 15828 15750 15840 15802
rect 15892 15750 15904 15802
rect 15956 15750 15968 15802
rect 16020 15750 16032 15802
rect 16084 15750 18860 15802
rect 1104 15728 18860 15750
rect 18138 15688 18144 15700
rect 18099 15660 18144 15688
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 1104 15258 18860 15280
rect 1104 15206 6880 15258
rect 6932 15206 6944 15258
rect 6996 15206 7008 15258
rect 7060 15206 7072 15258
rect 7124 15206 7136 15258
rect 7188 15206 12811 15258
rect 12863 15206 12875 15258
rect 12927 15206 12939 15258
rect 12991 15206 13003 15258
rect 13055 15206 13067 15258
rect 13119 15206 18860 15258
rect 1104 15184 18860 15206
rect 1104 14714 18860 14736
rect 1104 14662 3915 14714
rect 3967 14662 3979 14714
rect 4031 14662 4043 14714
rect 4095 14662 4107 14714
rect 4159 14662 4171 14714
rect 4223 14662 9846 14714
rect 9898 14662 9910 14714
rect 9962 14662 9974 14714
rect 10026 14662 10038 14714
rect 10090 14662 10102 14714
rect 10154 14662 15776 14714
rect 15828 14662 15840 14714
rect 15892 14662 15904 14714
rect 15956 14662 15968 14714
rect 16020 14662 16032 14714
rect 16084 14662 18860 14714
rect 1104 14640 18860 14662
rect 1104 14170 18860 14192
rect 1104 14118 6880 14170
rect 6932 14118 6944 14170
rect 6996 14118 7008 14170
rect 7060 14118 7072 14170
rect 7124 14118 7136 14170
rect 7188 14118 12811 14170
rect 12863 14118 12875 14170
rect 12927 14118 12939 14170
rect 12991 14118 13003 14170
rect 13055 14118 13067 14170
rect 13119 14118 18860 14170
rect 1104 14096 18860 14118
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 8294 13920 8300 13932
rect 1719 13892 8300 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 1104 13626 18860 13648
rect 1104 13574 3915 13626
rect 3967 13574 3979 13626
rect 4031 13574 4043 13626
rect 4095 13574 4107 13626
rect 4159 13574 4171 13626
rect 4223 13574 9846 13626
rect 9898 13574 9910 13626
rect 9962 13574 9974 13626
rect 10026 13574 10038 13626
rect 10090 13574 10102 13626
rect 10154 13574 15776 13626
rect 15828 13574 15840 13626
rect 15892 13574 15904 13626
rect 15956 13574 15968 13626
rect 16020 13574 16032 13626
rect 16084 13574 18860 13626
rect 1104 13552 18860 13574
rect 1394 13512 1400 13524
rect 1355 13484 1400 13512
rect 1394 13472 1400 13484
rect 1452 13472 1458 13524
rect 1104 13082 18860 13104
rect 1104 13030 6880 13082
rect 6932 13030 6944 13082
rect 6996 13030 7008 13082
rect 7060 13030 7072 13082
rect 7124 13030 7136 13082
rect 7188 13030 12811 13082
rect 12863 13030 12875 13082
rect 12927 13030 12939 13082
rect 12991 13030 13003 13082
rect 13055 13030 13067 13082
rect 13119 13030 18860 13082
rect 1104 13008 18860 13030
rect 1104 12538 18860 12560
rect 1104 12486 3915 12538
rect 3967 12486 3979 12538
rect 4031 12486 4043 12538
rect 4095 12486 4107 12538
rect 4159 12486 4171 12538
rect 4223 12486 9846 12538
rect 9898 12486 9910 12538
rect 9962 12486 9974 12538
rect 10026 12486 10038 12538
rect 10090 12486 10102 12538
rect 10154 12486 15776 12538
rect 15828 12486 15840 12538
rect 15892 12486 15904 12538
rect 15956 12486 15968 12538
rect 16020 12486 16032 12538
rect 16084 12486 18860 12538
rect 1104 12464 18860 12486
rect 1104 11994 18860 12016
rect 1104 11942 6880 11994
rect 6932 11942 6944 11994
rect 6996 11942 7008 11994
rect 7060 11942 7072 11994
rect 7124 11942 7136 11994
rect 7188 11942 12811 11994
rect 12863 11942 12875 11994
rect 12927 11942 12939 11994
rect 12991 11942 13003 11994
rect 13055 11942 13067 11994
rect 13119 11942 18860 11994
rect 1104 11920 18860 11942
rect 1104 11450 18860 11472
rect 1104 11398 3915 11450
rect 3967 11398 3979 11450
rect 4031 11398 4043 11450
rect 4095 11398 4107 11450
rect 4159 11398 4171 11450
rect 4223 11398 9846 11450
rect 9898 11398 9910 11450
rect 9962 11398 9974 11450
rect 10026 11398 10038 11450
rect 10090 11398 10102 11450
rect 10154 11398 15776 11450
rect 15828 11398 15840 11450
rect 15892 11398 15904 11450
rect 15956 11398 15968 11450
rect 16020 11398 16032 11450
rect 16084 11398 18860 11450
rect 1104 11376 18860 11398
rect 1104 10906 18860 10928
rect 1104 10854 6880 10906
rect 6932 10854 6944 10906
rect 6996 10854 7008 10906
rect 7060 10854 7072 10906
rect 7124 10854 7136 10906
rect 7188 10854 12811 10906
rect 12863 10854 12875 10906
rect 12927 10854 12939 10906
rect 12991 10854 13003 10906
rect 13055 10854 13067 10906
rect 13119 10854 18860 10906
rect 1104 10832 18860 10854
rect 1104 10362 18860 10384
rect 1104 10310 3915 10362
rect 3967 10310 3979 10362
rect 4031 10310 4043 10362
rect 4095 10310 4107 10362
rect 4159 10310 4171 10362
rect 4223 10310 9846 10362
rect 9898 10310 9910 10362
rect 9962 10310 9974 10362
rect 10026 10310 10038 10362
rect 10090 10310 10102 10362
rect 10154 10310 15776 10362
rect 15828 10310 15840 10362
rect 15892 10310 15904 10362
rect 15956 10310 15968 10362
rect 16020 10310 16032 10362
rect 16084 10310 18860 10362
rect 1104 10288 18860 10310
rect 1104 9818 18860 9840
rect 1104 9766 6880 9818
rect 6932 9766 6944 9818
rect 6996 9766 7008 9818
rect 7060 9766 7072 9818
rect 7124 9766 7136 9818
rect 7188 9766 12811 9818
rect 12863 9766 12875 9818
rect 12927 9766 12939 9818
rect 12991 9766 13003 9818
rect 13055 9766 13067 9818
rect 13119 9766 18860 9818
rect 1104 9744 18860 9766
rect 17405 9571 17463 9577
rect 17405 9537 17417 9571
rect 17451 9568 17463 9571
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17451 9540 17877 9568
rect 17451 9537 17463 9540
rect 17405 9531 17463 9537
rect 17865 9537 17877 9540
rect 17911 9568 17923 9571
rect 17954 9568 17960 9580
rect 17911 9540 17960 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18046 9432 18052 9444
rect 18007 9404 18052 9432
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 1104 9274 18860 9296
rect 1104 9222 3915 9274
rect 3967 9222 3979 9274
rect 4031 9222 4043 9274
rect 4095 9222 4107 9274
rect 4159 9222 4171 9274
rect 4223 9222 9846 9274
rect 9898 9222 9910 9274
rect 9962 9222 9974 9274
rect 10026 9222 10038 9274
rect 10090 9222 10102 9274
rect 10154 9222 15776 9274
rect 15828 9222 15840 9274
rect 15892 9222 15904 9274
rect 15956 9222 15968 9274
rect 16020 9222 16032 9274
rect 16084 9222 18860 9274
rect 1104 9200 18860 9222
rect 1104 8730 18860 8752
rect 1104 8678 6880 8730
rect 6932 8678 6944 8730
rect 6996 8678 7008 8730
rect 7060 8678 7072 8730
rect 7124 8678 7136 8730
rect 7188 8678 12811 8730
rect 12863 8678 12875 8730
rect 12927 8678 12939 8730
rect 12991 8678 13003 8730
rect 13055 8678 13067 8730
rect 13119 8678 18860 8730
rect 1104 8656 18860 8678
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1857 8483 1915 8489
rect 1857 8480 1869 8483
rect 1636 8452 1869 8480
rect 1636 8440 1642 8452
rect 1857 8449 1869 8452
rect 1903 8449 1915 8483
rect 1857 8443 1915 8449
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 11330 8344 11336 8356
rect 2087 8316 11336 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 1104 8186 18860 8208
rect 1104 8134 3915 8186
rect 3967 8134 3979 8186
rect 4031 8134 4043 8186
rect 4095 8134 4107 8186
rect 4159 8134 4171 8186
rect 4223 8134 9846 8186
rect 9898 8134 9910 8186
rect 9962 8134 9974 8186
rect 10026 8134 10038 8186
rect 10090 8134 10102 8186
rect 10154 8134 15776 8186
rect 15828 8134 15840 8186
rect 15892 8134 15904 8186
rect 15956 8134 15968 8186
rect 16020 8134 16032 8186
rect 16084 8134 18860 8186
rect 1104 8112 18860 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 1104 7642 18860 7664
rect 1104 7590 6880 7642
rect 6932 7590 6944 7642
rect 6996 7590 7008 7642
rect 7060 7590 7072 7642
rect 7124 7590 7136 7642
rect 7188 7590 12811 7642
rect 12863 7590 12875 7642
rect 12927 7590 12939 7642
rect 12991 7590 13003 7642
rect 13055 7590 13067 7642
rect 13119 7590 18860 7642
rect 1104 7568 18860 7590
rect 1104 7098 18860 7120
rect 1104 7046 3915 7098
rect 3967 7046 3979 7098
rect 4031 7046 4043 7098
rect 4095 7046 4107 7098
rect 4159 7046 4171 7098
rect 4223 7046 9846 7098
rect 9898 7046 9910 7098
rect 9962 7046 9974 7098
rect 10026 7046 10038 7098
rect 10090 7046 10102 7098
rect 10154 7046 15776 7098
rect 15828 7046 15840 7098
rect 15892 7046 15904 7098
rect 15956 7046 15968 7098
rect 16020 7046 16032 7098
rect 16084 7046 18860 7098
rect 1104 7024 18860 7046
rect 1104 6554 18860 6576
rect 1104 6502 6880 6554
rect 6932 6502 6944 6554
rect 6996 6502 7008 6554
rect 7060 6502 7072 6554
rect 7124 6502 7136 6554
rect 7188 6502 12811 6554
rect 12863 6502 12875 6554
rect 12927 6502 12939 6554
rect 12991 6502 13003 6554
rect 13055 6502 13067 6554
rect 13119 6502 18860 6554
rect 1104 6480 18860 6502
rect 1104 6010 18860 6032
rect 1104 5958 3915 6010
rect 3967 5958 3979 6010
rect 4031 5958 4043 6010
rect 4095 5958 4107 6010
rect 4159 5958 4171 6010
rect 4223 5958 9846 6010
rect 9898 5958 9910 6010
rect 9962 5958 9974 6010
rect 10026 5958 10038 6010
rect 10090 5958 10102 6010
rect 10154 5958 15776 6010
rect 15828 5958 15840 6010
rect 15892 5958 15904 6010
rect 15956 5958 15968 6010
rect 16020 5958 16032 6010
rect 16084 5958 18860 6010
rect 1104 5936 18860 5958
rect 1104 5466 18860 5488
rect 1104 5414 6880 5466
rect 6932 5414 6944 5466
rect 6996 5414 7008 5466
rect 7060 5414 7072 5466
rect 7124 5414 7136 5466
rect 7188 5414 12811 5466
rect 12863 5414 12875 5466
rect 12927 5414 12939 5466
rect 12991 5414 13003 5466
rect 13055 5414 13067 5466
rect 13119 5414 18860 5466
rect 1104 5392 18860 5414
rect 1104 4922 18860 4944
rect 1104 4870 3915 4922
rect 3967 4870 3979 4922
rect 4031 4870 4043 4922
rect 4095 4870 4107 4922
rect 4159 4870 4171 4922
rect 4223 4870 9846 4922
rect 9898 4870 9910 4922
rect 9962 4870 9974 4922
rect 10026 4870 10038 4922
rect 10090 4870 10102 4922
rect 10154 4870 15776 4922
rect 15828 4870 15840 4922
rect 15892 4870 15904 4922
rect 15956 4870 15968 4922
rect 16020 4870 16032 4922
rect 16084 4870 18860 4922
rect 1104 4848 18860 4870
rect 1104 4378 18860 4400
rect 1104 4326 6880 4378
rect 6932 4326 6944 4378
rect 6996 4326 7008 4378
rect 7060 4326 7072 4378
rect 7124 4326 7136 4378
rect 7188 4326 12811 4378
rect 12863 4326 12875 4378
rect 12927 4326 12939 4378
rect 12991 4326 13003 4378
rect 13055 4326 13067 4378
rect 13119 4326 18860 4378
rect 1104 4304 18860 4326
rect 1104 3834 18860 3856
rect 1104 3782 3915 3834
rect 3967 3782 3979 3834
rect 4031 3782 4043 3834
rect 4095 3782 4107 3834
rect 4159 3782 4171 3834
rect 4223 3782 9846 3834
rect 9898 3782 9910 3834
rect 9962 3782 9974 3834
rect 10026 3782 10038 3834
rect 10090 3782 10102 3834
rect 10154 3782 15776 3834
rect 15828 3782 15840 3834
rect 15892 3782 15904 3834
rect 15956 3782 15968 3834
rect 16020 3782 16032 3834
rect 16084 3782 18860 3834
rect 1104 3760 18860 3782
rect 16114 3476 16120 3528
rect 16172 3516 16178 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 16172 3488 17877 3516
rect 16172 3476 16178 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 1104 3290 18860 3312
rect 1104 3238 6880 3290
rect 6932 3238 6944 3290
rect 6996 3238 7008 3290
rect 7060 3238 7072 3290
rect 7124 3238 7136 3290
rect 7188 3238 12811 3290
rect 12863 3238 12875 3290
rect 12927 3238 12939 3290
rect 12991 3238 13003 3290
rect 13055 3238 13067 3290
rect 13119 3238 18860 3290
rect 1104 3216 18860 3238
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 1688 2972 1716 3003
rect 2222 2972 2228 2984
rect 1688 2944 2228 2972
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 1486 2836 1492 2848
rect 1447 2808 1492 2836
rect 1486 2796 1492 2808
rect 1544 2796 1550 2848
rect 1104 2746 18860 2768
rect 1104 2694 3915 2746
rect 3967 2694 3979 2746
rect 4031 2694 4043 2746
rect 4095 2694 4107 2746
rect 4159 2694 4171 2746
rect 4223 2694 9846 2746
rect 9898 2694 9910 2746
rect 9962 2694 9974 2746
rect 10026 2694 10038 2746
rect 10090 2694 10102 2746
rect 10154 2694 15776 2746
rect 15828 2694 15840 2746
rect 15892 2694 15904 2746
rect 15956 2694 15968 2746
rect 16020 2694 16032 2746
rect 16084 2694 18860 2746
rect 1104 2672 18860 2694
rect 12710 2632 12716 2644
rect 12671 2604 12716 2632
rect 12710 2592 12716 2604
rect 12768 2592 12774 2644
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 15436 2604 17693 2632
rect 15436 2592 15442 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 17681 2595 17739 2601
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 14734 2564 14740 2576
rect 8435 2536 14740 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8404 2428 8432 2527
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 7883 2400 8432 2428
rect 12069 2431 12127 2437
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12434 2428 12440 2440
rect 12115 2400 12440 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12434 2388 12440 2400
rect 12492 2428 12498 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12492 2400 12541 2428
rect 12492 2388 12498 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 17402 2428 17408 2440
rect 17083 2400 17408 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17402 2388 17408 2400
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 2133 2363 2191 2369
rect 2133 2329 2145 2363
rect 2179 2360 2191 2363
rect 2498 2360 2504 2372
rect 2179 2332 2504 2360
rect 2179 2329 2191 2332
rect 2133 2323 2191 2329
rect 2498 2320 2504 2332
rect 2556 2360 2562 2372
rect 2685 2363 2743 2369
rect 2685 2360 2697 2363
rect 2556 2332 2697 2360
rect 2556 2320 2562 2332
rect 2685 2329 2697 2332
rect 2731 2329 2743 2363
rect 2685 2323 2743 2329
rect 3053 2363 3111 2369
rect 3053 2329 3065 2363
rect 3099 2360 3111 2363
rect 13354 2360 13360 2372
rect 3099 2332 13360 2360
rect 3099 2329 3111 2332
rect 3053 2323 3111 2329
rect 13354 2320 13360 2332
rect 13412 2320 13418 2372
rect 7466 2252 7472 2304
rect 7524 2292 7530 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7524 2264 7665 2292
rect 7524 2252 7530 2264
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 1104 2202 18860 2224
rect 1104 2150 6880 2202
rect 6932 2150 6944 2202
rect 6996 2150 7008 2202
rect 7060 2150 7072 2202
rect 7124 2150 7136 2202
rect 7188 2150 12811 2202
rect 12863 2150 12875 2202
rect 12927 2150 12939 2202
rect 12991 2150 13003 2202
rect 13055 2150 13067 2202
rect 13119 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 18236 47404 18288 47456
rect 18420 47404 18472 47456
rect 3915 47302 3967 47354
rect 3979 47302 4031 47354
rect 4043 47302 4095 47354
rect 4107 47302 4159 47354
rect 4171 47302 4223 47354
rect 9846 47302 9898 47354
rect 9910 47302 9962 47354
rect 9974 47302 10026 47354
rect 10038 47302 10090 47354
rect 10102 47302 10154 47354
rect 15776 47302 15828 47354
rect 15840 47302 15892 47354
rect 15904 47302 15956 47354
rect 15968 47302 16020 47354
rect 16032 47302 16084 47354
rect 1492 47243 1544 47252
rect 1492 47209 1501 47243
rect 1501 47209 1535 47243
rect 1535 47209 1544 47243
rect 1492 47200 1544 47209
rect 10232 47243 10284 47252
rect 10232 47209 10241 47243
rect 10241 47209 10275 47243
rect 10275 47209 10284 47243
rect 10232 47200 10284 47209
rect 11060 47200 11112 47252
rect 11704 47200 11756 47252
rect 12440 47200 12492 47252
rect 14004 47132 14056 47184
rect 1124 47064 1176 47116
rect 2964 47064 3016 47116
rect 4252 47064 4304 47116
rect 4712 47064 4764 47116
rect 5724 47064 5776 47116
rect 7104 47064 7156 47116
rect 8944 47064 8996 47116
rect 16120 47107 16172 47116
rect 16120 47073 16129 47107
rect 16129 47073 16163 47107
rect 16163 47073 16172 47107
rect 16120 47064 16172 47073
rect 16488 47064 16540 47116
rect 1676 47039 1728 47048
rect 1676 47005 1685 47039
rect 1685 47005 1719 47039
rect 1719 47005 1728 47039
rect 1676 46996 1728 47005
rect 14832 47039 14884 47048
rect 14832 47005 14841 47039
rect 14841 47005 14875 47039
rect 14875 47005 14884 47039
rect 14832 46996 14884 47005
rect 15292 46996 15344 47048
rect 16856 46996 16908 47048
rect 2320 46860 2372 46912
rect 6184 46860 6236 46912
rect 8024 46860 8076 46912
rect 6880 46758 6932 46810
rect 6944 46758 6996 46810
rect 7008 46758 7060 46810
rect 7072 46758 7124 46810
rect 7136 46758 7188 46810
rect 12811 46758 12863 46810
rect 12875 46758 12927 46810
rect 12939 46758 12991 46810
rect 13003 46758 13055 46810
rect 13067 46758 13119 46810
rect 664 46656 716 46708
rect 1584 46656 1636 46708
rect 2688 46699 2740 46708
rect 2688 46665 2697 46699
rect 2697 46665 2731 46699
rect 2731 46665 2740 46699
rect 2688 46656 2740 46665
rect 3516 46699 3568 46708
rect 3516 46665 3525 46699
rect 3525 46665 3559 46699
rect 3559 46665 3568 46699
rect 3516 46656 3568 46665
rect 4896 46699 4948 46708
rect 4896 46665 4905 46699
rect 4905 46665 4939 46699
rect 4939 46665 4948 46699
rect 4896 46656 4948 46665
rect 5264 46656 5316 46708
rect 6736 46699 6788 46708
rect 6736 46665 6745 46699
rect 6745 46665 6779 46699
rect 6779 46665 6788 46699
rect 6736 46656 6788 46665
rect 7656 46699 7708 46708
rect 7656 46665 7665 46699
rect 7665 46665 7699 46699
rect 7699 46665 7708 46699
rect 7656 46656 7708 46665
rect 8576 46699 8628 46708
rect 8576 46665 8585 46699
rect 8585 46665 8619 46699
rect 8619 46665 8628 46699
rect 8576 46656 8628 46665
rect 14188 46699 14240 46708
rect 14188 46665 14197 46699
rect 14197 46665 14231 46699
rect 14231 46665 14240 46699
rect 14188 46656 14240 46665
rect 15476 46588 15528 46640
rect 16120 46656 16172 46708
rect 19156 46588 19208 46640
rect 9496 46563 9548 46572
rect 9496 46529 9505 46563
rect 9505 46529 9539 46563
rect 9539 46529 9548 46563
rect 9496 46520 9548 46529
rect 10508 46563 10560 46572
rect 10508 46529 10517 46563
rect 10517 46529 10551 46563
rect 10551 46529 10560 46563
rect 10508 46520 10560 46529
rect 11888 46563 11940 46572
rect 11888 46529 11897 46563
rect 11897 46529 11931 46563
rect 11931 46529 11940 46563
rect 11888 46520 11940 46529
rect 12716 46520 12768 46572
rect 13452 46563 13504 46572
rect 13452 46529 13461 46563
rect 13461 46529 13495 46563
rect 13495 46529 13504 46563
rect 13452 46520 13504 46529
rect 15108 46563 15160 46572
rect 15108 46529 15117 46563
rect 15117 46529 15151 46563
rect 15151 46529 15160 46563
rect 15108 46520 15160 46529
rect 15660 46520 15712 46572
rect 17316 46495 17368 46504
rect 17316 46461 17325 46495
rect 17325 46461 17359 46495
rect 17359 46461 17368 46495
rect 17316 46452 17368 46461
rect 19616 46452 19668 46504
rect 15568 46427 15620 46436
rect 15568 46393 15577 46427
rect 15577 46393 15611 46427
rect 15611 46393 15620 46427
rect 15568 46384 15620 46393
rect 3915 46214 3967 46266
rect 3979 46214 4031 46266
rect 4043 46214 4095 46266
rect 4107 46214 4159 46266
rect 4171 46214 4223 46266
rect 9846 46214 9898 46266
rect 9910 46214 9962 46266
rect 9974 46214 10026 46266
rect 10038 46214 10090 46266
rect 10102 46214 10154 46266
rect 15776 46214 15828 46266
rect 15840 46214 15892 46266
rect 15904 46214 15956 46266
rect 15968 46214 16020 46266
rect 16032 46214 16084 46266
rect 1676 46112 1728 46164
rect 2044 46155 2096 46164
rect 2044 46121 2053 46155
rect 2053 46121 2087 46155
rect 2087 46121 2096 46155
rect 2044 46112 2096 46121
rect 13636 46112 13688 46164
rect 14740 46155 14792 46164
rect 14740 46121 14749 46155
rect 14749 46121 14783 46155
rect 14783 46121 14792 46155
rect 14740 46112 14792 46121
rect 15476 46155 15528 46164
rect 15476 46121 15485 46155
rect 15485 46121 15519 46155
rect 15519 46121 15528 46155
rect 15476 46112 15528 46121
rect 17776 46112 17828 46164
rect 204 45976 256 46028
rect 16948 46019 17000 46028
rect 16948 45985 16957 46019
rect 16957 45985 16991 46019
rect 16991 45985 17000 46019
rect 16948 45976 17000 45985
rect 17040 45908 17092 45960
rect 17224 45951 17276 45960
rect 17224 45917 17233 45951
rect 17233 45917 17267 45951
rect 17267 45917 17276 45951
rect 17224 45908 17276 45917
rect 6880 45670 6932 45722
rect 6944 45670 6996 45722
rect 7008 45670 7060 45722
rect 7072 45670 7124 45722
rect 7136 45670 7188 45722
rect 12811 45670 12863 45722
rect 12875 45670 12927 45722
rect 12939 45670 12991 45722
rect 13003 45670 13055 45722
rect 13067 45670 13119 45722
rect 17316 45500 17368 45552
rect 17132 45475 17184 45484
rect 17132 45441 17141 45475
rect 17141 45441 17175 45475
rect 17175 45441 17184 45475
rect 17132 45432 17184 45441
rect 18052 45475 18104 45484
rect 18052 45441 18061 45475
rect 18061 45441 18095 45475
rect 18095 45441 18104 45475
rect 18052 45432 18104 45441
rect 18328 45432 18380 45484
rect 17408 45296 17460 45348
rect 17592 45296 17644 45348
rect 3915 45126 3967 45178
rect 3979 45126 4031 45178
rect 4043 45126 4095 45178
rect 4107 45126 4159 45178
rect 4171 45126 4223 45178
rect 9846 45126 9898 45178
rect 9910 45126 9962 45178
rect 9974 45126 10026 45178
rect 10038 45126 10090 45178
rect 10102 45126 10154 45178
rect 15776 45126 15828 45178
rect 15840 45126 15892 45178
rect 15904 45126 15956 45178
rect 15968 45126 16020 45178
rect 16032 45126 16084 45178
rect 16948 45024 17000 45076
rect 18052 45024 18104 45076
rect 18236 44820 18288 44872
rect 15476 44752 15528 44804
rect 6880 44582 6932 44634
rect 6944 44582 6996 44634
rect 7008 44582 7060 44634
rect 7072 44582 7124 44634
rect 7136 44582 7188 44634
rect 12811 44582 12863 44634
rect 12875 44582 12927 44634
rect 12939 44582 12991 44634
rect 13003 44582 13055 44634
rect 13067 44582 13119 44634
rect 16488 44480 16540 44532
rect 18236 44412 18288 44464
rect 18052 44344 18104 44396
rect 3915 44038 3967 44090
rect 3979 44038 4031 44090
rect 4043 44038 4095 44090
rect 4107 44038 4159 44090
rect 4171 44038 4223 44090
rect 9846 44038 9898 44090
rect 9910 44038 9962 44090
rect 9974 44038 10026 44090
rect 10038 44038 10090 44090
rect 10102 44038 10154 44090
rect 15776 44038 15828 44090
rect 15840 44038 15892 44090
rect 15904 44038 15956 44090
rect 15968 44038 16020 44090
rect 16032 44038 16084 44090
rect 6880 43494 6932 43546
rect 6944 43494 6996 43546
rect 7008 43494 7060 43546
rect 7072 43494 7124 43546
rect 7136 43494 7188 43546
rect 12811 43494 12863 43546
rect 12875 43494 12927 43546
rect 12939 43494 12991 43546
rect 13003 43494 13055 43546
rect 13067 43494 13119 43546
rect 3915 42950 3967 43002
rect 3979 42950 4031 43002
rect 4043 42950 4095 43002
rect 4107 42950 4159 43002
rect 4171 42950 4223 43002
rect 9846 42950 9898 43002
rect 9910 42950 9962 43002
rect 9974 42950 10026 43002
rect 10038 42950 10090 43002
rect 10102 42950 10154 43002
rect 15776 42950 15828 43002
rect 15840 42950 15892 43002
rect 15904 42950 15956 43002
rect 15968 42950 16020 43002
rect 16032 42950 16084 43002
rect 6880 42406 6932 42458
rect 6944 42406 6996 42458
rect 7008 42406 7060 42458
rect 7072 42406 7124 42458
rect 7136 42406 7188 42458
rect 12811 42406 12863 42458
rect 12875 42406 12927 42458
rect 12939 42406 12991 42458
rect 13003 42406 13055 42458
rect 13067 42406 13119 42458
rect 1676 42211 1728 42220
rect 1676 42177 1685 42211
rect 1685 42177 1719 42211
rect 1719 42177 1728 42211
rect 1676 42168 1728 42177
rect 1492 42007 1544 42016
rect 1492 41973 1501 42007
rect 1501 41973 1535 42007
rect 1535 41973 1544 42007
rect 1492 41964 1544 41973
rect 3915 41862 3967 41914
rect 3979 41862 4031 41914
rect 4043 41862 4095 41914
rect 4107 41862 4159 41914
rect 4171 41862 4223 41914
rect 9846 41862 9898 41914
rect 9910 41862 9962 41914
rect 9974 41862 10026 41914
rect 10038 41862 10090 41914
rect 10102 41862 10154 41914
rect 15776 41862 15828 41914
rect 15840 41862 15892 41914
rect 15904 41862 15956 41914
rect 15968 41862 16020 41914
rect 16032 41862 16084 41914
rect 6880 41318 6932 41370
rect 6944 41318 6996 41370
rect 7008 41318 7060 41370
rect 7072 41318 7124 41370
rect 7136 41318 7188 41370
rect 12811 41318 12863 41370
rect 12875 41318 12927 41370
rect 12939 41318 12991 41370
rect 13003 41318 13055 41370
rect 13067 41318 13119 41370
rect 18144 41123 18196 41132
rect 18144 41089 18153 41123
rect 18153 41089 18187 41123
rect 18187 41089 18196 41123
rect 18144 41080 18196 41089
rect 17960 40919 18012 40928
rect 17960 40885 17969 40919
rect 17969 40885 18003 40919
rect 18003 40885 18012 40919
rect 17960 40876 18012 40885
rect 3915 40774 3967 40826
rect 3979 40774 4031 40826
rect 4043 40774 4095 40826
rect 4107 40774 4159 40826
rect 4171 40774 4223 40826
rect 9846 40774 9898 40826
rect 9910 40774 9962 40826
rect 9974 40774 10026 40826
rect 10038 40774 10090 40826
rect 10102 40774 10154 40826
rect 15776 40774 15828 40826
rect 15840 40774 15892 40826
rect 15904 40774 15956 40826
rect 15968 40774 16020 40826
rect 16032 40774 16084 40826
rect 6880 40230 6932 40282
rect 6944 40230 6996 40282
rect 7008 40230 7060 40282
rect 7072 40230 7124 40282
rect 7136 40230 7188 40282
rect 12811 40230 12863 40282
rect 12875 40230 12927 40282
rect 12939 40230 12991 40282
rect 13003 40230 13055 40282
rect 13067 40230 13119 40282
rect 3915 39686 3967 39738
rect 3979 39686 4031 39738
rect 4043 39686 4095 39738
rect 4107 39686 4159 39738
rect 4171 39686 4223 39738
rect 9846 39686 9898 39738
rect 9910 39686 9962 39738
rect 9974 39686 10026 39738
rect 10038 39686 10090 39738
rect 10102 39686 10154 39738
rect 15776 39686 15828 39738
rect 15840 39686 15892 39738
rect 15904 39686 15956 39738
rect 15968 39686 16020 39738
rect 16032 39686 16084 39738
rect 6880 39142 6932 39194
rect 6944 39142 6996 39194
rect 7008 39142 7060 39194
rect 7072 39142 7124 39194
rect 7136 39142 7188 39194
rect 12811 39142 12863 39194
rect 12875 39142 12927 39194
rect 12939 39142 12991 39194
rect 13003 39142 13055 39194
rect 13067 39142 13119 39194
rect 3915 38598 3967 38650
rect 3979 38598 4031 38650
rect 4043 38598 4095 38650
rect 4107 38598 4159 38650
rect 4171 38598 4223 38650
rect 9846 38598 9898 38650
rect 9910 38598 9962 38650
rect 9974 38598 10026 38650
rect 10038 38598 10090 38650
rect 10102 38598 10154 38650
rect 15776 38598 15828 38650
rect 15840 38598 15892 38650
rect 15904 38598 15956 38650
rect 15968 38598 16020 38650
rect 16032 38598 16084 38650
rect 6880 38054 6932 38106
rect 6944 38054 6996 38106
rect 7008 38054 7060 38106
rect 7072 38054 7124 38106
rect 7136 38054 7188 38106
rect 12811 38054 12863 38106
rect 12875 38054 12927 38106
rect 12939 38054 12991 38106
rect 13003 38054 13055 38106
rect 13067 38054 13119 38106
rect 3915 37510 3967 37562
rect 3979 37510 4031 37562
rect 4043 37510 4095 37562
rect 4107 37510 4159 37562
rect 4171 37510 4223 37562
rect 9846 37510 9898 37562
rect 9910 37510 9962 37562
rect 9974 37510 10026 37562
rect 10038 37510 10090 37562
rect 10102 37510 10154 37562
rect 15776 37510 15828 37562
rect 15840 37510 15892 37562
rect 15904 37510 15956 37562
rect 15968 37510 16020 37562
rect 16032 37510 16084 37562
rect 17960 37247 18012 37256
rect 17960 37213 17969 37247
rect 17969 37213 18003 37247
rect 18003 37213 18012 37247
rect 17960 37204 18012 37213
rect 18144 37247 18196 37256
rect 18144 37213 18153 37247
rect 18153 37213 18187 37247
rect 18187 37213 18196 37247
rect 18144 37204 18196 37213
rect 16396 37136 16448 37188
rect 16948 37068 17000 37120
rect 6880 36966 6932 37018
rect 6944 36966 6996 37018
rect 7008 36966 7060 37018
rect 7072 36966 7124 37018
rect 7136 36966 7188 37018
rect 12811 36966 12863 37018
rect 12875 36966 12927 37018
rect 12939 36966 12991 37018
rect 13003 36966 13055 37018
rect 13067 36966 13119 37018
rect 17040 36864 17092 36916
rect 17960 36839 18012 36848
rect 17960 36805 17969 36839
rect 17969 36805 18003 36839
rect 18003 36805 18012 36839
rect 17960 36796 18012 36805
rect 18144 36771 18196 36780
rect 18144 36737 18153 36771
rect 18153 36737 18187 36771
rect 18187 36737 18196 36771
rect 18144 36728 18196 36737
rect 18236 36660 18288 36712
rect 17776 36567 17828 36576
rect 17776 36533 17785 36567
rect 17785 36533 17819 36567
rect 17819 36533 17828 36567
rect 17776 36524 17828 36533
rect 3915 36422 3967 36474
rect 3979 36422 4031 36474
rect 4043 36422 4095 36474
rect 4107 36422 4159 36474
rect 4171 36422 4223 36474
rect 9846 36422 9898 36474
rect 9910 36422 9962 36474
rect 9974 36422 10026 36474
rect 10038 36422 10090 36474
rect 10102 36422 10154 36474
rect 15776 36422 15828 36474
rect 15840 36422 15892 36474
rect 15904 36422 15956 36474
rect 15968 36422 16020 36474
rect 16032 36422 16084 36474
rect 18052 36363 18104 36372
rect 18052 36329 18061 36363
rect 18061 36329 18095 36363
rect 18095 36329 18104 36363
rect 18052 36320 18104 36329
rect 15200 36184 15252 36236
rect 16856 36116 16908 36168
rect 17960 36116 18012 36168
rect 1860 36091 1912 36100
rect 1860 36057 1869 36091
rect 1869 36057 1903 36091
rect 1903 36057 1912 36091
rect 1860 36048 1912 36057
rect 16580 36048 16632 36100
rect 17224 36048 17276 36100
rect 14280 35980 14332 36032
rect 15660 36023 15712 36032
rect 15660 35989 15669 36023
rect 15669 35989 15703 36023
rect 15703 35989 15712 36023
rect 15660 35980 15712 35989
rect 16304 36023 16356 36032
rect 16304 35989 16313 36023
rect 16313 35989 16347 36023
rect 16347 35989 16356 36023
rect 16304 35980 16356 35989
rect 6880 35878 6932 35930
rect 6944 35878 6996 35930
rect 7008 35878 7060 35930
rect 7072 35878 7124 35930
rect 7136 35878 7188 35930
rect 12811 35878 12863 35930
rect 12875 35878 12927 35930
rect 12939 35878 12991 35930
rect 13003 35878 13055 35930
rect 13067 35878 13119 35930
rect 1860 35776 1912 35828
rect 18144 35776 18196 35828
rect 15568 35708 15620 35760
rect 15660 35640 15712 35692
rect 16580 35640 16632 35692
rect 16856 35683 16908 35692
rect 16856 35649 16865 35683
rect 16865 35649 16899 35683
rect 16899 35649 16908 35683
rect 16856 35640 16908 35649
rect 17040 35640 17092 35692
rect 16212 35572 16264 35624
rect 18052 35572 18104 35624
rect 15108 35504 15160 35556
rect 14464 35436 14516 35488
rect 16856 35436 16908 35488
rect 3915 35334 3967 35386
rect 3979 35334 4031 35386
rect 4043 35334 4095 35386
rect 4107 35334 4159 35386
rect 4171 35334 4223 35386
rect 9846 35334 9898 35386
rect 9910 35334 9962 35386
rect 9974 35334 10026 35386
rect 10038 35334 10090 35386
rect 10102 35334 10154 35386
rect 15776 35334 15828 35386
rect 15840 35334 15892 35386
rect 15904 35334 15956 35386
rect 15968 35334 16020 35386
rect 16032 35334 16084 35386
rect 14372 35164 14424 35216
rect 16028 35164 16080 35216
rect 14832 35096 14884 35148
rect 17500 35232 17552 35284
rect 1676 35028 1728 35080
rect 15108 35028 15160 35080
rect 16580 35071 16632 35080
rect 2044 34960 2096 35012
rect 14924 34960 14976 35012
rect 16580 35037 16589 35071
rect 16589 35037 16623 35071
rect 16623 35037 16632 35071
rect 16580 35028 16632 35037
rect 17868 35028 17920 35080
rect 18144 34960 18196 35012
rect 16028 34892 16080 34944
rect 17776 34892 17828 34944
rect 6880 34790 6932 34842
rect 6944 34790 6996 34842
rect 7008 34790 7060 34842
rect 7072 34790 7124 34842
rect 7136 34790 7188 34842
rect 12811 34790 12863 34842
rect 12875 34790 12927 34842
rect 12939 34790 12991 34842
rect 13003 34790 13055 34842
rect 13067 34790 13119 34842
rect 15200 34688 15252 34740
rect 15476 34688 15528 34740
rect 14464 34620 14516 34672
rect 17960 34620 18012 34672
rect 14372 34552 14424 34604
rect 14740 34595 14792 34604
rect 14740 34561 14749 34595
rect 14749 34561 14783 34595
rect 14783 34561 14792 34595
rect 14740 34552 14792 34561
rect 14924 34595 14976 34604
rect 14924 34561 14933 34595
rect 14933 34561 14967 34595
rect 14967 34561 14976 34595
rect 14924 34552 14976 34561
rect 15016 34552 15068 34604
rect 13636 34459 13688 34468
rect 13636 34425 13645 34459
rect 13645 34425 13679 34459
rect 13679 34425 13688 34459
rect 13636 34416 13688 34425
rect 14832 34459 14884 34468
rect 14832 34425 14841 34459
rect 14841 34425 14875 34459
rect 14875 34425 14884 34459
rect 14832 34416 14884 34425
rect 15384 34484 15436 34536
rect 16396 34552 16448 34604
rect 16764 34552 16816 34604
rect 16948 34595 17000 34604
rect 16948 34561 16957 34595
rect 16957 34561 16991 34595
rect 16991 34561 17000 34595
rect 16948 34552 17000 34561
rect 16488 34484 16540 34536
rect 17868 34527 17920 34536
rect 17868 34493 17877 34527
rect 17877 34493 17911 34527
rect 17911 34493 17920 34527
rect 17868 34484 17920 34493
rect 17132 34416 17184 34468
rect 13452 34348 13504 34400
rect 16580 34348 16632 34400
rect 16948 34348 17000 34400
rect 3915 34246 3967 34298
rect 3979 34246 4031 34298
rect 4043 34246 4095 34298
rect 4107 34246 4159 34298
rect 4171 34246 4223 34298
rect 9846 34246 9898 34298
rect 9910 34246 9962 34298
rect 9974 34246 10026 34298
rect 10038 34246 10090 34298
rect 10102 34246 10154 34298
rect 15776 34246 15828 34298
rect 15840 34246 15892 34298
rect 15904 34246 15956 34298
rect 15968 34246 16020 34298
rect 16032 34246 16084 34298
rect 13452 34187 13504 34196
rect 13452 34153 13461 34187
rect 13461 34153 13495 34187
rect 13495 34153 13504 34187
rect 13452 34144 13504 34153
rect 16488 34144 16540 34196
rect 18052 34187 18104 34196
rect 18052 34153 18061 34187
rect 18061 34153 18095 34187
rect 18095 34153 18104 34187
rect 18052 34144 18104 34153
rect 13636 34008 13688 34060
rect 15660 34008 15712 34060
rect 16396 34051 16448 34060
rect 14464 33940 14516 33992
rect 15476 33983 15528 33992
rect 15476 33949 15485 33983
rect 15485 33949 15519 33983
rect 15519 33949 15528 33983
rect 15476 33940 15528 33949
rect 16028 33940 16080 33992
rect 16396 34017 16405 34051
rect 16405 34017 16439 34051
rect 16439 34017 16448 34051
rect 16396 34008 16448 34017
rect 17960 34076 18012 34128
rect 17500 34008 17552 34060
rect 17684 34008 17736 34060
rect 18144 34051 18196 34060
rect 16672 33940 16724 33992
rect 17040 33940 17092 33992
rect 17776 33940 17828 33992
rect 18144 34017 18153 34051
rect 18153 34017 18187 34051
rect 18187 34017 18196 34051
rect 18144 34008 18196 34017
rect 14648 33915 14700 33924
rect 14648 33881 14657 33915
rect 14657 33881 14691 33915
rect 14691 33881 14700 33915
rect 14648 33872 14700 33881
rect 15568 33872 15620 33924
rect 12716 33847 12768 33856
rect 12716 33813 12725 33847
rect 12725 33813 12759 33847
rect 12759 33813 12768 33847
rect 12716 33804 12768 33813
rect 13452 33804 13504 33856
rect 14924 33804 14976 33856
rect 15108 33804 15160 33856
rect 16580 33872 16632 33924
rect 6880 33702 6932 33754
rect 6944 33702 6996 33754
rect 7008 33702 7060 33754
rect 7072 33702 7124 33754
rect 7136 33702 7188 33754
rect 12811 33702 12863 33754
rect 12875 33702 12927 33754
rect 12939 33702 12991 33754
rect 13003 33702 13055 33754
rect 13067 33702 13119 33754
rect 14740 33600 14792 33652
rect 14924 33600 14976 33652
rect 14280 33575 14332 33584
rect 13452 33507 13504 33516
rect 13452 33473 13461 33507
rect 13461 33473 13495 33507
rect 13495 33473 13504 33507
rect 13452 33464 13504 33473
rect 13544 33464 13596 33516
rect 14280 33541 14289 33575
rect 14289 33541 14323 33575
rect 14323 33541 14332 33575
rect 14280 33532 14332 33541
rect 15200 33532 15252 33584
rect 14556 33464 14608 33516
rect 14648 33464 14700 33516
rect 15568 33600 15620 33652
rect 15016 33396 15068 33448
rect 16028 33532 16080 33584
rect 16764 33532 16816 33584
rect 15844 33507 15896 33516
rect 15844 33473 15853 33507
rect 15853 33473 15887 33507
rect 15887 33473 15896 33507
rect 16948 33507 17000 33516
rect 15844 33464 15896 33473
rect 16948 33473 16957 33507
rect 16957 33473 16991 33507
rect 16991 33473 17000 33507
rect 16948 33464 17000 33473
rect 17408 33507 17460 33516
rect 17408 33473 17417 33507
rect 17417 33473 17451 33507
rect 17451 33473 17460 33507
rect 17408 33464 17460 33473
rect 17960 33464 18012 33516
rect 16212 33396 16264 33448
rect 17500 33439 17552 33448
rect 17500 33405 17509 33439
rect 17509 33405 17543 33439
rect 17543 33405 17552 33439
rect 17500 33396 17552 33405
rect 16856 33328 16908 33380
rect 17868 33328 17920 33380
rect 14740 33260 14792 33312
rect 15200 33260 15252 33312
rect 16304 33260 16356 33312
rect 3915 33158 3967 33210
rect 3979 33158 4031 33210
rect 4043 33158 4095 33210
rect 4107 33158 4159 33210
rect 4171 33158 4223 33210
rect 9846 33158 9898 33210
rect 9910 33158 9962 33210
rect 9974 33158 10026 33210
rect 10038 33158 10090 33210
rect 10102 33158 10154 33210
rect 15776 33158 15828 33210
rect 15840 33158 15892 33210
rect 15904 33158 15956 33210
rect 15968 33158 16020 33210
rect 16032 33158 16084 33210
rect 15108 33099 15160 33108
rect 15108 33065 15117 33099
rect 15117 33065 15151 33099
rect 15151 33065 15160 33099
rect 15108 33056 15160 33065
rect 14740 32988 14792 33040
rect 14556 32920 14608 32972
rect 14280 32895 14332 32904
rect 14280 32861 14289 32895
rect 14289 32861 14323 32895
rect 14323 32861 14332 32895
rect 14280 32852 14332 32861
rect 15200 32852 15252 32904
rect 16304 32895 16356 32904
rect 12716 32716 12768 32768
rect 13360 32716 13412 32768
rect 14832 32784 14884 32836
rect 16304 32861 16313 32895
rect 16313 32861 16347 32895
rect 16347 32861 16356 32895
rect 16304 32852 16356 32861
rect 16580 33056 16632 33108
rect 16856 33056 16908 33108
rect 17500 32920 17552 32972
rect 17776 32920 17828 32972
rect 16856 32895 16908 32904
rect 16856 32861 16865 32895
rect 16865 32861 16899 32895
rect 16899 32861 16908 32895
rect 16856 32852 16908 32861
rect 16948 32852 17000 32904
rect 17040 32716 17092 32768
rect 17316 32716 17368 32768
rect 6880 32614 6932 32666
rect 6944 32614 6996 32666
rect 7008 32614 7060 32666
rect 7072 32614 7124 32666
rect 7136 32614 7188 32666
rect 12811 32614 12863 32666
rect 12875 32614 12927 32666
rect 12939 32614 12991 32666
rect 13003 32614 13055 32666
rect 13067 32614 13119 32666
rect 13636 32555 13688 32564
rect 13636 32521 13645 32555
rect 13645 32521 13679 32555
rect 13679 32521 13688 32555
rect 13636 32512 13688 32521
rect 15200 32512 15252 32564
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 15292 32444 15344 32496
rect 16948 32512 17000 32564
rect 17408 32555 17460 32564
rect 17408 32521 17417 32555
rect 17417 32521 17451 32555
rect 17451 32521 17460 32555
rect 17408 32512 17460 32521
rect 18144 32512 18196 32564
rect 14740 32419 14792 32428
rect 14740 32385 14749 32419
rect 14749 32385 14783 32419
rect 14783 32385 14792 32419
rect 14740 32376 14792 32385
rect 14832 32419 14884 32428
rect 14832 32385 14841 32419
rect 14841 32385 14875 32419
rect 14875 32385 14884 32419
rect 14832 32376 14884 32385
rect 15568 32376 15620 32428
rect 16580 32376 16632 32428
rect 17592 32444 17644 32496
rect 16764 32376 16816 32428
rect 16856 32419 16908 32428
rect 16856 32385 16865 32419
rect 16865 32385 16899 32419
rect 16899 32385 16908 32419
rect 16856 32376 16908 32385
rect 17040 32376 17092 32428
rect 15016 32172 15068 32224
rect 15200 32215 15252 32224
rect 15200 32181 15209 32215
rect 15209 32181 15243 32215
rect 15243 32181 15252 32215
rect 15200 32172 15252 32181
rect 16028 32240 16080 32292
rect 16672 32240 16724 32292
rect 17132 32240 17184 32292
rect 17684 32240 17736 32292
rect 16580 32172 16632 32224
rect 3915 32070 3967 32122
rect 3979 32070 4031 32122
rect 4043 32070 4095 32122
rect 4107 32070 4159 32122
rect 4171 32070 4223 32122
rect 9846 32070 9898 32122
rect 9910 32070 9962 32122
rect 9974 32070 10026 32122
rect 10038 32070 10090 32122
rect 10102 32070 10154 32122
rect 15776 32070 15828 32122
rect 15840 32070 15892 32122
rect 15904 32070 15956 32122
rect 15968 32070 16020 32122
rect 16032 32070 16084 32122
rect 15016 31968 15068 32020
rect 15476 31968 15528 32020
rect 17040 31968 17092 32020
rect 17500 31968 17552 32020
rect 14740 31875 14792 31884
rect 14740 31841 14749 31875
rect 14749 31841 14783 31875
rect 14783 31841 14792 31875
rect 14740 31832 14792 31841
rect 13360 31764 13412 31816
rect 17684 31900 17736 31952
rect 16856 31832 16908 31884
rect 16764 31764 16816 31816
rect 17316 31764 17368 31816
rect 17500 31764 17552 31816
rect 17408 31696 17460 31748
rect 6880 31526 6932 31578
rect 6944 31526 6996 31578
rect 7008 31526 7060 31578
rect 7072 31526 7124 31578
rect 7136 31526 7188 31578
rect 12811 31526 12863 31578
rect 12875 31526 12927 31578
rect 12939 31526 12991 31578
rect 13003 31526 13055 31578
rect 13067 31526 13119 31578
rect 15568 31424 15620 31476
rect 17040 31424 17092 31476
rect 17960 31467 18012 31476
rect 17960 31433 17969 31467
rect 17969 31433 18003 31467
rect 18003 31433 18012 31467
rect 17960 31424 18012 31433
rect 12716 31356 12768 31408
rect 16580 31356 16632 31408
rect 14096 31288 14148 31340
rect 16488 31288 16540 31340
rect 16948 31288 17000 31340
rect 17132 31331 17184 31340
rect 17132 31297 17141 31331
rect 17141 31297 17175 31331
rect 17175 31297 17184 31331
rect 17132 31288 17184 31297
rect 17684 31331 17736 31340
rect 17684 31297 17693 31331
rect 17693 31297 17727 31331
rect 17727 31297 17736 31331
rect 17684 31288 17736 31297
rect 15292 31220 15344 31272
rect 16120 31152 16172 31204
rect 16672 31084 16724 31136
rect 3915 30982 3967 31034
rect 3979 30982 4031 31034
rect 4043 30982 4095 31034
rect 4107 30982 4159 31034
rect 4171 30982 4223 31034
rect 9846 30982 9898 31034
rect 9910 30982 9962 31034
rect 9974 30982 10026 31034
rect 10038 30982 10090 31034
rect 10102 30982 10154 31034
rect 15776 30982 15828 31034
rect 15840 30982 15892 31034
rect 15904 30982 15956 31034
rect 15968 30982 16020 31034
rect 16032 30982 16084 31034
rect 17408 30923 17460 30932
rect 17408 30889 17417 30923
rect 17417 30889 17451 30923
rect 17451 30889 17460 30923
rect 17408 30880 17460 30889
rect 15200 30812 15252 30864
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 14096 30676 14148 30728
rect 15476 30676 15528 30728
rect 16028 30719 16080 30728
rect 16028 30685 16037 30719
rect 16037 30685 16071 30719
rect 16071 30685 16080 30719
rect 16028 30676 16080 30685
rect 18144 30812 18196 30864
rect 17776 30744 17828 30796
rect 17500 30719 17552 30728
rect 17500 30685 17509 30719
rect 17509 30685 17543 30719
rect 17543 30685 17552 30719
rect 17500 30676 17552 30685
rect 15752 30540 15804 30592
rect 6880 30438 6932 30490
rect 6944 30438 6996 30490
rect 7008 30438 7060 30490
rect 7072 30438 7124 30490
rect 7136 30438 7188 30490
rect 12811 30438 12863 30490
rect 12875 30438 12927 30490
rect 12939 30438 12991 30490
rect 13003 30438 13055 30490
rect 13067 30438 13119 30490
rect 1400 30379 1452 30388
rect 1400 30345 1409 30379
rect 1409 30345 1443 30379
rect 1443 30345 1452 30379
rect 1400 30336 1452 30345
rect 17316 30379 17368 30388
rect 17316 30345 17325 30379
rect 17325 30345 17359 30379
rect 17359 30345 17368 30379
rect 17316 30336 17368 30345
rect 15384 30268 15436 30320
rect 15752 30243 15804 30252
rect 15752 30209 15761 30243
rect 15761 30209 15795 30243
rect 15795 30209 15804 30243
rect 15752 30200 15804 30209
rect 15108 30132 15160 30184
rect 16028 30200 16080 30252
rect 17132 30200 17184 30252
rect 17868 30200 17920 30252
rect 18052 30200 18104 30252
rect 17592 30064 17644 30116
rect 3915 29894 3967 29946
rect 3979 29894 4031 29946
rect 4043 29894 4095 29946
rect 4107 29894 4159 29946
rect 4171 29894 4223 29946
rect 9846 29894 9898 29946
rect 9910 29894 9962 29946
rect 9974 29894 10026 29946
rect 10038 29894 10090 29946
rect 10102 29894 10154 29946
rect 15776 29894 15828 29946
rect 15840 29894 15892 29946
rect 15904 29894 15956 29946
rect 15968 29894 16020 29946
rect 16032 29894 16084 29946
rect 14372 29656 14424 29708
rect 15108 29656 15160 29708
rect 15660 29588 15712 29640
rect 17132 29588 17184 29640
rect 13636 29452 13688 29504
rect 15568 29452 15620 29504
rect 17960 29452 18012 29504
rect 6880 29350 6932 29402
rect 6944 29350 6996 29402
rect 7008 29350 7060 29402
rect 7072 29350 7124 29402
rect 7136 29350 7188 29402
rect 12811 29350 12863 29402
rect 12875 29350 12927 29402
rect 12939 29350 12991 29402
rect 13003 29350 13055 29402
rect 13067 29350 13119 29402
rect 3915 28806 3967 28858
rect 3979 28806 4031 28858
rect 4043 28806 4095 28858
rect 4107 28806 4159 28858
rect 4171 28806 4223 28858
rect 9846 28806 9898 28858
rect 9910 28806 9962 28858
rect 9974 28806 10026 28858
rect 10038 28806 10090 28858
rect 10102 28806 10154 28858
rect 15776 28806 15828 28858
rect 15840 28806 15892 28858
rect 15904 28806 15956 28858
rect 15968 28806 16020 28858
rect 16032 28806 16084 28858
rect 16212 28704 16264 28756
rect 18144 28543 18196 28552
rect 18144 28509 18153 28543
rect 18153 28509 18187 28543
rect 18187 28509 18196 28543
rect 18144 28500 18196 28509
rect 6880 28262 6932 28314
rect 6944 28262 6996 28314
rect 7008 28262 7060 28314
rect 7072 28262 7124 28314
rect 7136 28262 7188 28314
rect 12811 28262 12863 28314
rect 12875 28262 12927 28314
rect 12939 28262 12991 28314
rect 13003 28262 13055 28314
rect 13067 28262 13119 28314
rect 3915 27718 3967 27770
rect 3979 27718 4031 27770
rect 4043 27718 4095 27770
rect 4107 27718 4159 27770
rect 4171 27718 4223 27770
rect 9846 27718 9898 27770
rect 9910 27718 9962 27770
rect 9974 27718 10026 27770
rect 10038 27718 10090 27770
rect 10102 27718 10154 27770
rect 15776 27718 15828 27770
rect 15840 27718 15892 27770
rect 15904 27718 15956 27770
rect 15968 27718 16020 27770
rect 16032 27718 16084 27770
rect 6880 27174 6932 27226
rect 6944 27174 6996 27226
rect 7008 27174 7060 27226
rect 7072 27174 7124 27226
rect 7136 27174 7188 27226
rect 12811 27174 12863 27226
rect 12875 27174 12927 27226
rect 12939 27174 12991 27226
rect 13003 27174 13055 27226
rect 13067 27174 13119 27226
rect 3915 26630 3967 26682
rect 3979 26630 4031 26682
rect 4043 26630 4095 26682
rect 4107 26630 4159 26682
rect 4171 26630 4223 26682
rect 9846 26630 9898 26682
rect 9910 26630 9962 26682
rect 9974 26630 10026 26682
rect 10038 26630 10090 26682
rect 10102 26630 10154 26682
rect 15776 26630 15828 26682
rect 15840 26630 15892 26682
rect 15904 26630 15956 26682
rect 15968 26630 16020 26682
rect 16032 26630 16084 26682
rect 6880 26086 6932 26138
rect 6944 26086 6996 26138
rect 7008 26086 7060 26138
rect 7072 26086 7124 26138
rect 7136 26086 7188 26138
rect 12811 26086 12863 26138
rect 12875 26086 12927 26138
rect 12939 26086 12991 26138
rect 13003 26086 13055 26138
rect 13067 26086 13119 26138
rect 14372 26027 14424 26036
rect 14372 25993 14381 26027
rect 14381 25993 14415 26027
rect 14415 25993 14424 26027
rect 14372 25984 14424 25993
rect 13636 25848 13688 25900
rect 13452 25780 13504 25832
rect 14188 25823 14240 25832
rect 14188 25789 14197 25823
rect 14197 25789 14231 25823
rect 14231 25789 14240 25823
rect 14188 25780 14240 25789
rect 3915 25542 3967 25594
rect 3979 25542 4031 25594
rect 4043 25542 4095 25594
rect 4107 25542 4159 25594
rect 4171 25542 4223 25594
rect 9846 25542 9898 25594
rect 9910 25542 9962 25594
rect 9974 25542 10026 25594
rect 10038 25542 10090 25594
rect 10102 25542 10154 25594
rect 15776 25542 15828 25594
rect 15840 25542 15892 25594
rect 15904 25542 15956 25594
rect 15968 25542 16020 25594
rect 16032 25542 16084 25594
rect 13176 25483 13228 25492
rect 13176 25449 13185 25483
rect 13185 25449 13219 25483
rect 13219 25449 13228 25483
rect 13176 25440 13228 25449
rect 11152 25236 11204 25288
rect 1492 25143 1544 25152
rect 1492 25109 1501 25143
rect 1501 25109 1535 25143
rect 1535 25109 1544 25143
rect 1492 25100 1544 25109
rect 6880 24998 6932 25050
rect 6944 24998 6996 25050
rect 7008 24998 7060 25050
rect 7072 24998 7124 25050
rect 7136 24998 7188 25050
rect 12811 24998 12863 25050
rect 12875 24998 12927 25050
rect 12939 24998 12991 25050
rect 13003 24998 13055 25050
rect 13067 24998 13119 25050
rect 13176 24828 13228 24880
rect 1676 24760 1728 24812
rect 12532 24760 12584 24812
rect 13452 24803 13504 24812
rect 13452 24769 13461 24803
rect 13461 24769 13495 24803
rect 13495 24769 13504 24803
rect 13452 24760 13504 24769
rect 14188 24760 14240 24812
rect 13544 24599 13596 24608
rect 13544 24565 13553 24599
rect 13553 24565 13587 24599
rect 13587 24565 13596 24599
rect 13544 24556 13596 24565
rect 3915 24454 3967 24506
rect 3979 24454 4031 24506
rect 4043 24454 4095 24506
rect 4107 24454 4159 24506
rect 4171 24454 4223 24506
rect 9846 24454 9898 24506
rect 9910 24454 9962 24506
rect 9974 24454 10026 24506
rect 10038 24454 10090 24506
rect 10102 24454 10154 24506
rect 15776 24454 15828 24506
rect 15840 24454 15892 24506
rect 15904 24454 15956 24506
rect 15968 24454 16020 24506
rect 16032 24454 16084 24506
rect 13452 24352 13504 24404
rect 11152 24327 11204 24336
rect 11152 24293 11161 24327
rect 11161 24293 11195 24327
rect 11195 24293 11204 24327
rect 11152 24284 11204 24293
rect 13176 24327 13228 24336
rect 13176 24293 13185 24327
rect 13185 24293 13219 24327
rect 13219 24293 13228 24327
rect 13176 24284 13228 24293
rect 13544 24216 13596 24268
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 13176 24148 13228 24200
rect 13636 24080 13688 24132
rect 6880 23910 6932 23962
rect 6944 23910 6996 23962
rect 7008 23910 7060 23962
rect 7072 23910 7124 23962
rect 7136 23910 7188 23962
rect 12811 23910 12863 23962
rect 12875 23910 12927 23962
rect 12939 23910 12991 23962
rect 13003 23910 13055 23962
rect 13067 23910 13119 23962
rect 3915 23366 3967 23418
rect 3979 23366 4031 23418
rect 4043 23366 4095 23418
rect 4107 23366 4159 23418
rect 4171 23366 4223 23418
rect 9846 23366 9898 23418
rect 9910 23366 9962 23418
rect 9974 23366 10026 23418
rect 10038 23366 10090 23418
rect 10102 23366 10154 23418
rect 15776 23366 15828 23418
rect 15840 23366 15892 23418
rect 15904 23366 15956 23418
rect 15968 23366 16020 23418
rect 16032 23366 16084 23418
rect 6880 22822 6932 22874
rect 6944 22822 6996 22874
rect 7008 22822 7060 22874
rect 7072 22822 7124 22874
rect 7136 22822 7188 22874
rect 12811 22822 12863 22874
rect 12875 22822 12927 22874
rect 12939 22822 12991 22874
rect 13003 22822 13055 22874
rect 13067 22822 13119 22874
rect 3915 22278 3967 22330
rect 3979 22278 4031 22330
rect 4043 22278 4095 22330
rect 4107 22278 4159 22330
rect 4171 22278 4223 22330
rect 9846 22278 9898 22330
rect 9910 22278 9962 22330
rect 9974 22278 10026 22330
rect 10038 22278 10090 22330
rect 10102 22278 10154 22330
rect 15776 22278 15828 22330
rect 15840 22278 15892 22330
rect 15904 22278 15956 22330
rect 15968 22278 16020 22330
rect 16032 22278 16084 22330
rect 13636 22040 13688 22092
rect 14004 22040 14056 22092
rect 13452 21972 13504 22024
rect 18144 22015 18196 22024
rect 18144 21981 18153 22015
rect 18153 21981 18187 22015
rect 18187 21981 18196 22015
rect 18144 21972 18196 21981
rect 13268 21836 13320 21888
rect 18052 21836 18104 21888
rect 6880 21734 6932 21786
rect 6944 21734 6996 21786
rect 7008 21734 7060 21786
rect 7072 21734 7124 21786
rect 7136 21734 7188 21786
rect 12811 21734 12863 21786
rect 12875 21734 12927 21786
rect 12939 21734 12991 21786
rect 13003 21734 13055 21786
rect 13067 21734 13119 21786
rect 3915 21190 3967 21242
rect 3979 21190 4031 21242
rect 4043 21190 4095 21242
rect 4107 21190 4159 21242
rect 4171 21190 4223 21242
rect 9846 21190 9898 21242
rect 9910 21190 9962 21242
rect 9974 21190 10026 21242
rect 10038 21190 10090 21242
rect 10102 21190 10154 21242
rect 15776 21190 15828 21242
rect 15840 21190 15892 21242
rect 15904 21190 15956 21242
rect 15968 21190 16020 21242
rect 16032 21190 16084 21242
rect 6880 20646 6932 20698
rect 6944 20646 6996 20698
rect 7008 20646 7060 20698
rect 7072 20646 7124 20698
rect 7136 20646 7188 20698
rect 12811 20646 12863 20698
rect 12875 20646 12927 20698
rect 12939 20646 12991 20698
rect 13003 20646 13055 20698
rect 13067 20646 13119 20698
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 15016 20204 15068 20256
rect 3915 20102 3967 20154
rect 3979 20102 4031 20154
rect 4043 20102 4095 20154
rect 4107 20102 4159 20154
rect 4171 20102 4223 20154
rect 9846 20102 9898 20154
rect 9910 20102 9962 20154
rect 9974 20102 10026 20154
rect 10038 20102 10090 20154
rect 10102 20102 10154 20154
rect 15776 20102 15828 20154
rect 15840 20102 15892 20154
rect 15904 20102 15956 20154
rect 15968 20102 16020 20154
rect 16032 20102 16084 20154
rect 1676 19907 1728 19916
rect 1676 19873 1685 19907
rect 1685 19873 1719 19907
rect 1719 19873 1728 19907
rect 1676 19864 1728 19873
rect 1400 19839 1452 19848
rect 1400 19805 1409 19839
rect 1409 19805 1443 19839
rect 1443 19805 1452 19839
rect 1400 19796 1452 19805
rect 6880 19558 6932 19610
rect 6944 19558 6996 19610
rect 7008 19558 7060 19610
rect 7072 19558 7124 19610
rect 7136 19558 7188 19610
rect 12811 19558 12863 19610
rect 12875 19558 12927 19610
rect 12939 19558 12991 19610
rect 13003 19558 13055 19610
rect 13067 19558 13119 19610
rect 1400 19431 1452 19440
rect 1400 19397 1409 19431
rect 1409 19397 1443 19431
rect 1443 19397 1452 19431
rect 1400 19388 1452 19397
rect 14004 19252 14056 19304
rect 15016 19252 15068 19304
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 3915 19014 3967 19066
rect 3979 19014 4031 19066
rect 4043 19014 4095 19066
rect 4107 19014 4159 19066
rect 4171 19014 4223 19066
rect 9846 19014 9898 19066
rect 9910 19014 9962 19066
rect 9974 19014 10026 19066
rect 10038 19014 10090 19066
rect 10102 19014 10154 19066
rect 15776 19014 15828 19066
rect 15840 19014 15892 19066
rect 15904 19014 15956 19066
rect 15968 19014 16020 19066
rect 16032 19014 16084 19066
rect 6880 18470 6932 18522
rect 6944 18470 6996 18522
rect 7008 18470 7060 18522
rect 7072 18470 7124 18522
rect 7136 18470 7188 18522
rect 12811 18470 12863 18522
rect 12875 18470 12927 18522
rect 12939 18470 12991 18522
rect 13003 18470 13055 18522
rect 13067 18470 13119 18522
rect 13452 18368 13504 18420
rect 13268 18300 13320 18352
rect 8300 18164 8352 18216
rect 11336 18232 11388 18284
rect 3915 17926 3967 17978
rect 3979 17926 4031 17978
rect 4043 17926 4095 17978
rect 4107 17926 4159 17978
rect 4171 17926 4223 17978
rect 9846 17926 9898 17978
rect 9910 17926 9962 17978
rect 9974 17926 10026 17978
rect 10038 17926 10090 17978
rect 10102 17926 10154 17978
rect 15776 17926 15828 17978
rect 15840 17926 15892 17978
rect 15904 17926 15956 17978
rect 15968 17926 16020 17978
rect 16032 17926 16084 17978
rect 11336 17527 11388 17536
rect 11336 17493 11345 17527
rect 11345 17493 11379 17527
rect 11379 17493 11388 17527
rect 11336 17484 11388 17493
rect 6880 17382 6932 17434
rect 6944 17382 6996 17434
rect 7008 17382 7060 17434
rect 7072 17382 7124 17434
rect 7136 17382 7188 17434
rect 12811 17382 12863 17434
rect 12875 17382 12927 17434
rect 12939 17382 12991 17434
rect 13003 17382 13055 17434
rect 13067 17382 13119 17434
rect 3915 16838 3967 16890
rect 3979 16838 4031 16890
rect 4043 16838 4095 16890
rect 4107 16838 4159 16890
rect 4171 16838 4223 16890
rect 9846 16838 9898 16890
rect 9910 16838 9962 16890
rect 9974 16838 10026 16890
rect 10038 16838 10090 16890
rect 10102 16838 10154 16890
rect 15776 16838 15828 16890
rect 15840 16838 15892 16890
rect 15904 16838 15956 16890
rect 15968 16838 16020 16890
rect 16032 16838 16084 16890
rect 6880 16294 6932 16346
rect 6944 16294 6996 16346
rect 7008 16294 7060 16346
rect 7072 16294 7124 16346
rect 7136 16294 7188 16346
rect 12811 16294 12863 16346
rect 12875 16294 12927 16346
rect 12939 16294 12991 16346
rect 13003 16294 13055 16346
rect 13067 16294 13119 16346
rect 17868 16099 17920 16108
rect 17868 16065 17877 16099
rect 17877 16065 17911 16099
rect 17911 16065 17920 16099
rect 17868 16056 17920 16065
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 3915 15750 3967 15802
rect 3979 15750 4031 15802
rect 4043 15750 4095 15802
rect 4107 15750 4159 15802
rect 4171 15750 4223 15802
rect 9846 15750 9898 15802
rect 9910 15750 9962 15802
rect 9974 15750 10026 15802
rect 10038 15750 10090 15802
rect 10102 15750 10154 15802
rect 15776 15750 15828 15802
rect 15840 15750 15892 15802
rect 15904 15750 15956 15802
rect 15968 15750 16020 15802
rect 16032 15750 16084 15802
rect 18144 15691 18196 15700
rect 18144 15657 18153 15691
rect 18153 15657 18187 15691
rect 18187 15657 18196 15691
rect 18144 15648 18196 15657
rect 6880 15206 6932 15258
rect 6944 15206 6996 15258
rect 7008 15206 7060 15258
rect 7072 15206 7124 15258
rect 7136 15206 7188 15258
rect 12811 15206 12863 15258
rect 12875 15206 12927 15258
rect 12939 15206 12991 15258
rect 13003 15206 13055 15258
rect 13067 15206 13119 15258
rect 3915 14662 3967 14714
rect 3979 14662 4031 14714
rect 4043 14662 4095 14714
rect 4107 14662 4159 14714
rect 4171 14662 4223 14714
rect 9846 14662 9898 14714
rect 9910 14662 9962 14714
rect 9974 14662 10026 14714
rect 10038 14662 10090 14714
rect 10102 14662 10154 14714
rect 15776 14662 15828 14714
rect 15840 14662 15892 14714
rect 15904 14662 15956 14714
rect 15968 14662 16020 14714
rect 16032 14662 16084 14714
rect 6880 14118 6932 14170
rect 6944 14118 6996 14170
rect 7008 14118 7060 14170
rect 7072 14118 7124 14170
rect 7136 14118 7188 14170
rect 12811 14118 12863 14170
rect 12875 14118 12927 14170
rect 12939 14118 12991 14170
rect 13003 14118 13055 14170
rect 13067 14118 13119 14170
rect 8300 13880 8352 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 3915 13574 3967 13626
rect 3979 13574 4031 13626
rect 4043 13574 4095 13626
rect 4107 13574 4159 13626
rect 4171 13574 4223 13626
rect 9846 13574 9898 13626
rect 9910 13574 9962 13626
rect 9974 13574 10026 13626
rect 10038 13574 10090 13626
rect 10102 13574 10154 13626
rect 15776 13574 15828 13626
rect 15840 13574 15892 13626
rect 15904 13574 15956 13626
rect 15968 13574 16020 13626
rect 16032 13574 16084 13626
rect 1400 13515 1452 13524
rect 1400 13481 1409 13515
rect 1409 13481 1443 13515
rect 1443 13481 1452 13515
rect 1400 13472 1452 13481
rect 6880 13030 6932 13082
rect 6944 13030 6996 13082
rect 7008 13030 7060 13082
rect 7072 13030 7124 13082
rect 7136 13030 7188 13082
rect 12811 13030 12863 13082
rect 12875 13030 12927 13082
rect 12939 13030 12991 13082
rect 13003 13030 13055 13082
rect 13067 13030 13119 13082
rect 3915 12486 3967 12538
rect 3979 12486 4031 12538
rect 4043 12486 4095 12538
rect 4107 12486 4159 12538
rect 4171 12486 4223 12538
rect 9846 12486 9898 12538
rect 9910 12486 9962 12538
rect 9974 12486 10026 12538
rect 10038 12486 10090 12538
rect 10102 12486 10154 12538
rect 15776 12486 15828 12538
rect 15840 12486 15892 12538
rect 15904 12486 15956 12538
rect 15968 12486 16020 12538
rect 16032 12486 16084 12538
rect 6880 11942 6932 11994
rect 6944 11942 6996 11994
rect 7008 11942 7060 11994
rect 7072 11942 7124 11994
rect 7136 11942 7188 11994
rect 12811 11942 12863 11994
rect 12875 11942 12927 11994
rect 12939 11942 12991 11994
rect 13003 11942 13055 11994
rect 13067 11942 13119 11994
rect 3915 11398 3967 11450
rect 3979 11398 4031 11450
rect 4043 11398 4095 11450
rect 4107 11398 4159 11450
rect 4171 11398 4223 11450
rect 9846 11398 9898 11450
rect 9910 11398 9962 11450
rect 9974 11398 10026 11450
rect 10038 11398 10090 11450
rect 10102 11398 10154 11450
rect 15776 11398 15828 11450
rect 15840 11398 15892 11450
rect 15904 11398 15956 11450
rect 15968 11398 16020 11450
rect 16032 11398 16084 11450
rect 6880 10854 6932 10906
rect 6944 10854 6996 10906
rect 7008 10854 7060 10906
rect 7072 10854 7124 10906
rect 7136 10854 7188 10906
rect 12811 10854 12863 10906
rect 12875 10854 12927 10906
rect 12939 10854 12991 10906
rect 13003 10854 13055 10906
rect 13067 10854 13119 10906
rect 3915 10310 3967 10362
rect 3979 10310 4031 10362
rect 4043 10310 4095 10362
rect 4107 10310 4159 10362
rect 4171 10310 4223 10362
rect 9846 10310 9898 10362
rect 9910 10310 9962 10362
rect 9974 10310 10026 10362
rect 10038 10310 10090 10362
rect 10102 10310 10154 10362
rect 15776 10310 15828 10362
rect 15840 10310 15892 10362
rect 15904 10310 15956 10362
rect 15968 10310 16020 10362
rect 16032 10310 16084 10362
rect 6880 9766 6932 9818
rect 6944 9766 6996 9818
rect 7008 9766 7060 9818
rect 7072 9766 7124 9818
rect 7136 9766 7188 9818
rect 12811 9766 12863 9818
rect 12875 9766 12927 9818
rect 12939 9766 12991 9818
rect 13003 9766 13055 9818
rect 13067 9766 13119 9818
rect 17960 9528 18012 9580
rect 18052 9435 18104 9444
rect 18052 9401 18061 9435
rect 18061 9401 18095 9435
rect 18095 9401 18104 9435
rect 18052 9392 18104 9401
rect 3915 9222 3967 9274
rect 3979 9222 4031 9274
rect 4043 9222 4095 9274
rect 4107 9222 4159 9274
rect 4171 9222 4223 9274
rect 9846 9222 9898 9274
rect 9910 9222 9962 9274
rect 9974 9222 10026 9274
rect 10038 9222 10090 9274
rect 10102 9222 10154 9274
rect 15776 9222 15828 9274
rect 15840 9222 15892 9274
rect 15904 9222 15956 9274
rect 15968 9222 16020 9274
rect 16032 9222 16084 9274
rect 6880 8678 6932 8730
rect 6944 8678 6996 8730
rect 7008 8678 7060 8730
rect 7072 8678 7124 8730
rect 7136 8678 7188 8730
rect 12811 8678 12863 8730
rect 12875 8678 12927 8730
rect 12939 8678 12991 8730
rect 13003 8678 13055 8730
rect 13067 8678 13119 8730
rect 1584 8440 1636 8492
rect 11336 8304 11388 8356
rect 3915 8134 3967 8186
rect 3979 8134 4031 8186
rect 4043 8134 4095 8186
rect 4107 8134 4159 8186
rect 4171 8134 4223 8186
rect 9846 8134 9898 8186
rect 9910 8134 9962 8186
rect 9974 8134 10026 8186
rect 10038 8134 10090 8186
rect 10102 8134 10154 8186
rect 15776 8134 15828 8186
rect 15840 8134 15892 8186
rect 15904 8134 15956 8186
rect 15968 8134 16020 8186
rect 16032 8134 16084 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 6880 7590 6932 7642
rect 6944 7590 6996 7642
rect 7008 7590 7060 7642
rect 7072 7590 7124 7642
rect 7136 7590 7188 7642
rect 12811 7590 12863 7642
rect 12875 7590 12927 7642
rect 12939 7590 12991 7642
rect 13003 7590 13055 7642
rect 13067 7590 13119 7642
rect 3915 7046 3967 7098
rect 3979 7046 4031 7098
rect 4043 7046 4095 7098
rect 4107 7046 4159 7098
rect 4171 7046 4223 7098
rect 9846 7046 9898 7098
rect 9910 7046 9962 7098
rect 9974 7046 10026 7098
rect 10038 7046 10090 7098
rect 10102 7046 10154 7098
rect 15776 7046 15828 7098
rect 15840 7046 15892 7098
rect 15904 7046 15956 7098
rect 15968 7046 16020 7098
rect 16032 7046 16084 7098
rect 6880 6502 6932 6554
rect 6944 6502 6996 6554
rect 7008 6502 7060 6554
rect 7072 6502 7124 6554
rect 7136 6502 7188 6554
rect 12811 6502 12863 6554
rect 12875 6502 12927 6554
rect 12939 6502 12991 6554
rect 13003 6502 13055 6554
rect 13067 6502 13119 6554
rect 3915 5958 3967 6010
rect 3979 5958 4031 6010
rect 4043 5958 4095 6010
rect 4107 5958 4159 6010
rect 4171 5958 4223 6010
rect 9846 5958 9898 6010
rect 9910 5958 9962 6010
rect 9974 5958 10026 6010
rect 10038 5958 10090 6010
rect 10102 5958 10154 6010
rect 15776 5958 15828 6010
rect 15840 5958 15892 6010
rect 15904 5958 15956 6010
rect 15968 5958 16020 6010
rect 16032 5958 16084 6010
rect 6880 5414 6932 5466
rect 6944 5414 6996 5466
rect 7008 5414 7060 5466
rect 7072 5414 7124 5466
rect 7136 5414 7188 5466
rect 12811 5414 12863 5466
rect 12875 5414 12927 5466
rect 12939 5414 12991 5466
rect 13003 5414 13055 5466
rect 13067 5414 13119 5466
rect 3915 4870 3967 4922
rect 3979 4870 4031 4922
rect 4043 4870 4095 4922
rect 4107 4870 4159 4922
rect 4171 4870 4223 4922
rect 9846 4870 9898 4922
rect 9910 4870 9962 4922
rect 9974 4870 10026 4922
rect 10038 4870 10090 4922
rect 10102 4870 10154 4922
rect 15776 4870 15828 4922
rect 15840 4870 15892 4922
rect 15904 4870 15956 4922
rect 15968 4870 16020 4922
rect 16032 4870 16084 4922
rect 6880 4326 6932 4378
rect 6944 4326 6996 4378
rect 7008 4326 7060 4378
rect 7072 4326 7124 4378
rect 7136 4326 7188 4378
rect 12811 4326 12863 4378
rect 12875 4326 12927 4378
rect 12939 4326 12991 4378
rect 13003 4326 13055 4378
rect 13067 4326 13119 4378
rect 3915 3782 3967 3834
rect 3979 3782 4031 3834
rect 4043 3782 4095 3834
rect 4107 3782 4159 3834
rect 4171 3782 4223 3834
rect 9846 3782 9898 3834
rect 9910 3782 9962 3834
rect 9974 3782 10026 3834
rect 10038 3782 10090 3834
rect 10102 3782 10154 3834
rect 15776 3782 15828 3834
rect 15840 3782 15892 3834
rect 15904 3782 15956 3834
rect 15968 3782 16020 3834
rect 16032 3782 16084 3834
rect 16120 3476 16172 3528
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 6880 3238 6932 3290
rect 6944 3238 6996 3290
rect 7008 3238 7060 3290
rect 7072 3238 7124 3290
rect 7136 3238 7188 3290
rect 12811 3238 12863 3290
rect 12875 3238 12927 3290
rect 12939 3238 12991 3290
rect 13003 3238 13055 3290
rect 13067 3238 13119 3290
rect 2228 2975 2280 2984
rect 2228 2941 2237 2975
rect 2237 2941 2271 2975
rect 2271 2941 2280 2975
rect 2228 2932 2280 2941
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 3915 2694 3967 2746
rect 3979 2694 4031 2746
rect 4043 2694 4095 2746
rect 4107 2694 4159 2746
rect 4171 2694 4223 2746
rect 9846 2694 9898 2746
rect 9910 2694 9962 2746
rect 9974 2694 10026 2746
rect 10038 2694 10090 2746
rect 10102 2694 10154 2746
rect 15776 2694 15828 2746
rect 15840 2694 15892 2746
rect 15904 2694 15956 2746
rect 15968 2694 16020 2746
rect 16032 2694 16084 2746
rect 12716 2635 12768 2644
rect 12716 2601 12725 2635
rect 12725 2601 12759 2635
rect 12759 2601 12768 2635
rect 12716 2592 12768 2601
rect 15384 2592 15436 2644
rect 14740 2524 14792 2576
rect 12440 2388 12492 2440
rect 17408 2388 17460 2440
rect 2504 2320 2556 2372
rect 13360 2320 13412 2372
rect 7472 2252 7524 2304
rect 6880 2150 6932 2202
rect 6944 2150 6996 2202
rect 7008 2150 7060 2202
rect 7072 2150 7124 2202
rect 7136 2150 7188 2202
rect 12811 2150 12863 2202
rect 12875 2150 12927 2202
rect 12939 2150 12991 2202
rect 13003 2150 13055 2202
rect 13067 2150 13119 2202
<< metal2 >>
rect 202 49200 258 50000
rect 662 49200 718 50000
rect 1122 49200 1178 50000
rect 1582 49200 1638 50000
rect 2042 49314 2098 50000
rect 2502 49314 2558 50000
rect 2042 49286 2360 49314
rect 2042 49200 2098 49286
rect 216 46034 244 49200
rect 676 46714 704 49200
rect 1136 47122 1164 49200
rect 1490 47288 1546 47297
rect 1490 47223 1492 47232
rect 1544 47223 1546 47232
rect 1492 47194 1544 47200
rect 1124 47116 1176 47122
rect 1124 47058 1176 47064
rect 1596 46714 1624 49200
rect 1676 47048 1728 47054
rect 1676 46990 1728 46996
rect 664 46708 716 46714
rect 664 46650 716 46656
rect 1584 46708 1636 46714
rect 1584 46650 1636 46656
rect 1688 46170 1716 46990
rect 2332 46918 2360 49286
rect 2502 49286 2728 49314
rect 2502 49200 2558 49286
rect 2320 46912 2372 46918
rect 2320 46854 2372 46860
rect 2700 46714 2728 49286
rect 2962 49200 3018 50000
rect 3422 49314 3478 50000
rect 3882 49314 3938 50000
rect 4342 49314 4398 50000
rect 4802 49314 4858 50000
rect 3422 49286 3556 49314
rect 3422 49200 3478 49286
rect 2976 47122 3004 49200
rect 2964 47116 3016 47122
rect 2964 47058 3016 47064
rect 3528 46714 3556 49286
rect 3882 49286 4108 49314
rect 3882 49200 3938 49286
rect 4080 47546 4108 49286
rect 4342 49286 4752 49314
rect 4342 49200 4398 49286
rect 4080 47518 4292 47546
rect 3915 47356 4223 47376
rect 3915 47354 3921 47356
rect 3977 47354 4001 47356
rect 4057 47354 4081 47356
rect 4137 47354 4161 47356
rect 4217 47354 4223 47356
rect 3977 47302 3979 47354
rect 4159 47302 4161 47354
rect 3915 47300 3921 47302
rect 3977 47300 4001 47302
rect 4057 47300 4081 47302
rect 4137 47300 4161 47302
rect 4217 47300 4223 47302
rect 3915 47280 4223 47300
rect 4264 47122 4292 47518
rect 4724 47122 4752 49286
rect 4802 49286 4936 49314
rect 4802 49200 4858 49286
rect 4252 47116 4304 47122
rect 4252 47058 4304 47064
rect 4712 47116 4764 47122
rect 4712 47058 4764 47064
rect 4908 46714 4936 49286
rect 5262 49200 5318 50000
rect 5722 49200 5778 50000
rect 6182 49200 6238 50000
rect 6642 49314 6698 50000
rect 6642 49286 6776 49314
rect 6642 49200 6698 49286
rect 5276 46714 5304 49200
rect 5736 47122 5764 49200
rect 5724 47116 5776 47122
rect 5724 47058 5776 47064
rect 6196 46918 6224 49200
rect 6184 46912 6236 46918
rect 6184 46854 6236 46860
rect 6748 46714 6776 49286
rect 7102 49200 7158 50000
rect 7562 49314 7618 50000
rect 7562 49286 7696 49314
rect 7562 49200 7618 49286
rect 7116 47122 7144 49200
rect 7104 47116 7156 47122
rect 7104 47058 7156 47064
rect 6880 46812 7188 46832
rect 6880 46810 6886 46812
rect 6942 46810 6966 46812
rect 7022 46810 7046 46812
rect 7102 46810 7126 46812
rect 7182 46810 7188 46812
rect 6942 46758 6944 46810
rect 7124 46758 7126 46810
rect 6880 46756 6886 46758
rect 6942 46756 6966 46758
rect 7022 46756 7046 46758
rect 7102 46756 7126 46758
rect 7182 46756 7188 46758
rect 6880 46736 7188 46756
rect 7668 46714 7696 49286
rect 8022 49200 8078 50000
rect 8482 49314 8538 50000
rect 8482 49286 8616 49314
rect 8482 49200 8538 49286
rect 8036 46918 8064 49200
rect 8024 46912 8076 46918
rect 8024 46854 8076 46860
rect 8588 46714 8616 49286
rect 8942 49200 8998 50000
rect 9402 49314 9458 50000
rect 9862 49314 9918 50000
rect 10414 49314 10470 50000
rect 10874 49314 10930 50000
rect 11334 49314 11390 50000
rect 11794 49314 11850 50000
rect 12254 49314 12310 50000
rect 9402 49286 9536 49314
rect 9402 49200 9458 49286
rect 8956 47122 8984 49200
rect 8944 47116 8996 47122
rect 8944 47058 8996 47064
rect 2688 46708 2740 46714
rect 2688 46650 2740 46656
rect 3516 46708 3568 46714
rect 3516 46650 3568 46656
rect 4896 46708 4948 46714
rect 4896 46650 4948 46656
rect 5264 46708 5316 46714
rect 5264 46650 5316 46656
rect 6736 46708 6788 46714
rect 6736 46650 6788 46656
rect 7656 46708 7708 46714
rect 7656 46650 7708 46656
rect 8576 46708 8628 46714
rect 8576 46650 8628 46656
rect 9508 46578 9536 49286
rect 9862 49286 10272 49314
rect 9862 49200 9918 49286
rect 9846 47356 10154 47376
rect 9846 47354 9852 47356
rect 9908 47354 9932 47356
rect 9988 47354 10012 47356
rect 10068 47354 10092 47356
rect 10148 47354 10154 47356
rect 9908 47302 9910 47354
rect 10090 47302 10092 47354
rect 9846 47300 9852 47302
rect 9908 47300 9932 47302
rect 9988 47300 10012 47302
rect 10068 47300 10092 47302
rect 10148 47300 10154 47302
rect 9846 47280 10154 47300
rect 10244 47258 10272 49286
rect 10414 49286 10548 49314
rect 10414 49200 10470 49286
rect 10232 47252 10284 47258
rect 10232 47194 10284 47200
rect 10520 46578 10548 49286
rect 10874 49286 11008 49314
rect 10874 49200 10930 49286
rect 10980 47274 11008 49286
rect 11334 49286 11744 49314
rect 11334 49200 11390 49286
rect 10980 47258 11100 47274
rect 11716 47258 11744 49286
rect 11794 49286 11928 49314
rect 11794 49200 11850 49286
rect 10980 47252 11112 47258
rect 10980 47246 11060 47252
rect 11060 47194 11112 47200
rect 11704 47252 11756 47258
rect 11704 47194 11756 47200
rect 11900 46578 11928 49286
rect 12254 49286 12388 49314
rect 12254 49200 12310 49286
rect 12360 47274 12388 49286
rect 12714 49200 12770 50000
rect 13174 49314 13230 50000
rect 13174 49286 13492 49314
rect 13174 49200 13230 49286
rect 12360 47258 12480 47274
rect 12360 47252 12492 47258
rect 12360 47246 12440 47252
rect 12440 47194 12492 47200
rect 12728 46578 12756 49200
rect 12811 46812 13119 46832
rect 12811 46810 12817 46812
rect 12873 46810 12897 46812
rect 12953 46810 12977 46812
rect 13033 46810 13057 46812
rect 13113 46810 13119 46812
rect 12873 46758 12875 46810
rect 13055 46758 13057 46810
rect 12811 46756 12817 46758
rect 12873 46756 12897 46758
rect 12953 46756 12977 46758
rect 13033 46756 13057 46758
rect 13113 46756 13119 46758
rect 12811 46736 13119 46756
rect 13464 46578 13492 49286
rect 13634 49200 13690 50000
rect 14094 49314 14150 50000
rect 14554 49314 14610 50000
rect 15014 49314 15070 50000
rect 14094 49286 14228 49314
rect 14094 49200 14150 49286
rect 9496 46572 9548 46578
rect 9496 46514 9548 46520
rect 10508 46572 10560 46578
rect 10508 46514 10560 46520
rect 11888 46572 11940 46578
rect 11888 46514 11940 46520
rect 12716 46572 12768 46578
rect 12716 46514 12768 46520
rect 13452 46572 13504 46578
rect 13452 46514 13504 46520
rect 3915 46268 4223 46288
rect 3915 46266 3921 46268
rect 3977 46266 4001 46268
rect 4057 46266 4081 46268
rect 4137 46266 4161 46268
rect 4217 46266 4223 46268
rect 3977 46214 3979 46266
rect 4159 46214 4161 46266
rect 3915 46212 3921 46214
rect 3977 46212 4001 46214
rect 4057 46212 4081 46214
rect 4137 46212 4161 46214
rect 4217 46212 4223 46214
rect 3915 46192 4223 46212
rect 9846 46268 10154 46288
rect 9846 46266 9852 46268
rect 9908 46266 9932 46268
rect 9988 46266 10012 46268
rect 10068 46266 10092 46268
rect 10148 46266 10154 46268
rect 9908 46214 9910 46266
rect 10090 46214 10092 46266
rect 9846 46212 9852 46214
rect 9908 46212 9932 46214
rect 9988 46212 10012 46214
rect 10068 46212 10092 46214
rect 10148 46212 10154 46214
rect 9846 46192 10154 46212
rect 13648 46170 13676 49200
rect 14004 47184 14056 47190
rect 14004 47126 14056 47132
rect 1676 46164 1728 46170
rect 1676 46106 1728 46112
rect 2044 46164 2096 46170
rect 2044 46106 2096 46112
rect 13636 46164 13688 46170
rect 13636 46106 13688 46112
rect 204 46028 256 46034
rect 204 45970 256 45976
rect 1676 42220 1728 42226
rect 1676 42162 1728 42168
rect 1492 42016 1544 42022
rect 1492 41958 1544 41964
rect 1504 41721 1532 41958
rect 1490 41712 1546 41721
rect 1490 41647 1546 41656
rect 1688 35086 1716 42162
rect 1858 36136 1914 36145
rect 1858 36071 1860 36080
rect 1912 36071 1914 36080
rect 1860 36042 1912 36048
rect 1872 35834 1900 36042
rect 1860 35828 1912 35834
rect 1860 35770 1912 35776
rect 1676 35080 1728 35086
rect 1676 35022 1728 35028
rect 2056 35018 2084 46106
rect 6880 45724 7188 45744
rect 6880 45722 6886 45724
rect 6942 45722 6966 45724
rect 7022 45722 7046 45724
rect 7102 45722 7126 45724
rect 7182 45722 7188 45724
rect 6942 45670 6944 45722
rect 7124 45670 7126 45722
rect 6880 45668 6886 45670
rect 6942 45668 6966 45670
rect 7022 45668 7046 45670
rect 7102 45668 7126 45670
rect 7182 45668 7188 45670
rect 6880 45648 7188 45668
rect 12811 45724 13119 45744
rect 12811 45722 12817 45724
rect 12873 45722 12897 45724
rect 12953 45722 12977 45724
rect 13033 45722 13057 45724
rect 13113 45722 13119 45724
rect 12873 45670 12875 45722
rect 13055 45670 13057 45722
rect 12811 45668 12817 45670
rect 12873 45668 12897 45670
rect 12953 45668 12977 45670
rect 13033 45668 13057 45670
rect 13113 45668 13119 45670
rect 12811 45648 13119 45668
rect 3915 45180 4223 45200
rect 3915 45178 3921 45180
rect 3977 45178 4001 45180
rect 4057 45178 4081 45180
rect 4137 45178 4161 45180
rect 4217 45178 4223 45180
rect 3977 45126 3979 45178
rect 4159 45126 4161 45178
rect 3915 45124 3921 45126
rect 3977 45124 4001 45126
rect 4057 45124 4081 45126
rect 4137 45124 4161 45126
rect 4217 45124 4223 45126
rect 3915 45104 4223 45124
rect 9846 45180 10154 45200
rect 9846 45178 9852 45180
rect 9908 45178 9932 45180
rect 9988 45178 10012 45180
rect 10068 45178 10092 45180
rect 10148 45178 10154 45180
rect 9908 45126 9910 45178
rect 10090 45126 10092 45178
rect 9846 45124 9852 45126
rect 9908 45124 9932 45126
rect 9988 45124 10012 45126
rect 10068 45124 10092 45126
rect 10148 45124 10154 45126
rect 9846 45104 10154 45124
rect 6880 44636 7188 44656
rect 6880 44634 6886 44636
rect 6942 44634 6966 44636
rect 7022 44634 7046 44636
rect 7102 44634 7126 44636
rect 7182 44634 7188 44636
rect 6942 44582 6944 44634
rect 7124 44582 7126 44634
rect 6880 44580 6886 44582
rect 6942 44580 6966 44582
rect 7022 44580 7046 44582
rect 7102 44580 7126 44582
rect 7182 44580 7188 44582
rect 6880 44560 7188 44580
rect 12811 44636 13119 44656
rect 12811 44634 12817 44636
rect 12873 44634 12897 44636
rect 12953 44634 12977 44636
rect 13033 44634 13057 44636
rect 13113 44634 13119 44636
rect 12873 44582 12875 44634
rect 13055 44582 13057 44634
rect 12811 44580 12817 44582
rect 12873 44580 12897 44582
rect 12953 44580 12977 44582
rect 13033 44580 13057 44582
rect 13113 44580 13119 44582
rect 12811 44560 13119 44580
rect 3915 44092 4223 44112
rect 3915 44090 3921 44092
rect 3977 44090 4001 44092
rect 4057 44090 4081 44092
rect 4137 44090 4161 44092
rect 4217 44090 4223 44092
rect 3977 44038 3979 44090
rect 4159 44038 4161 44090
rect 3915 44036 3921 44038
rect 3977 44036 4001 44038
rect 4057 44036 4081 44038
rect 4137 44036 4161 44038
rect 4217 44036 4223 44038
rect 3915 44016 4223 44036
rect 9846 44092 10154 44112
rect 9846 44090 9852 44092
rect 9908 44090 9932 44092
rect 9988 44090 10012 44092
rect 10068 44090 10092 44092
rect 10148 44090 10154 44092
rect 9908 44038 9910 44090
rect 10090 44038 10092 44090
rect 9846 44036 9852 44038
rect 9908 44036 9932 44038
rect 9988 44036 10012 44038
rect 10068 44036 10092 44038
rect 10148 44036 10154 44038
rect 9846 44016 10154 44036
rect 6880 43548 7188 43568
rect 6880 43546 6886 43548
rect 6942 43546 6966 43548
rect 7022 43546 7046 43548
rect 7102 43546 7126 43548
rect 7182 43546 7188 43548
rect 6942 43494 6944 43546
rect 7124 43494 7126 43546
rect 6880 43492 6886 43494
rect 6942 43492 6966 43494
rect 7022 43492 7046 43494
rect 7102 43492 7126 43494
rect 7182 43492 7188 43494
rect 6880 43472 7188 43492
rect 12811 43548 13119 43568
rect 12811 43546 12817 43548
rect 12873 43546 12897 43548
rect 12953 43546 12977 43548
rect 13033 43546 13057 43548
rect 13113 43546 13119 43548
rect 12873 43494 12875 43546
rect 13055 43494 13057 43546
rect 12811 43492 12817 43494
rect 12873 43492 12897 43494
rect 12953 43492 12977 43494
rect 13033 43492 13057 43494
rect 13113 43492 13119 43494
rect 12811 43472 13119 43492
rect 3915 43004 4223 43024
rect 3915 43002 3921 43004
rect 3977 43002 4001 43004
rect 4057 43002 4081 43004
rect 4137 43002 4161 43004
rect 4217 43002 4223 43004
rect 3977 42950 3979 43002
rect 4159 42950 4161 43002
rect 3915 42948 3921 42950
rect 3977 42948 4001 42950
rect 4057 42948 4081 42950
rect 4137 42948 4161 42950
rect 4217 42948 4223 42950
rect 3915 42928 4223 42948
rect 9846 43004 10154 43024
rect 9846 43002 9852 43004
rect 9908 43002 9932 43004
rect 9988 43002 10012 43004
rect 10068 43002 10092 43004
rect 10148 43002 10154 43004
rect 9908 42950 9910 43002
rect 10090 42950 10092 43002
rect 9846 42948 9852 42950
rect 9908 42948 9932 42950
rect 9988 42948 10012 42950
rect 10068 42948 10092 42950
rect 10148 42948 10154 42950
rect 9846 42928 10154 42948
rect 6880 42460 7188 42480
rect 6880 42458 6886 42460
rect 6942 42458 6966 42460
rect 7022 42458 7046 42460
rect 7102 42458 7126 42460
rect 7182 42458 7188 42460
rect 6942 42406 6944 42458
rect 7124 42406 7126 42458
rect 6880 42404 6886 42406
rect 6942 42404 6966 42406
rect 7022 42404 7046 42406
rect 7102 42404 7126 42406
rect 7182 42404 7188 42406
rect 6880 42384 7188 42404
rect 12811 42460 13119 42480
rect 12811 42458 12817 42460
rect 12873 42458 12897 42460
rect 12953 42458 12977 42460
rect 13033 42458 13057 42460
rect 13113 42458 13119 42460
rect 12873 42406 12875 42458
rect 13055 42406 13057 42458
rect 12811 42404 12817 42406
rect 12873 42404 12897 42406
rect 12953 42404 12977 42406
rect 13033 42404 13057 42406
rect 13113 42404 13119 42406
rect 12811 42384 13119 42404
rect 3915 41916 4223 41936
rect 3915 41914 3921 41916
rect 3977 41914 4001 41916
rect 4057 41914 4081 41916
rect 4137 41914 4161 41916
rect 4217 41914 4223 41916
rect 3977 41862 3979 41914
rect 4159 41862 4161 41914
rect 3915 41860 3921 41862
rect 3977 41860 4001 41862
rect 4057 41860 4081 41862
rect 4137 41860 4161 41862
rect 4217 41860 4223 41862
rect 3915 41840 4223 41860
rect 9846 41916 10154 41936
rect 9846 41914 9852 41916
rect 9908 41914 9932 41916
rect 9988 41914 10012 41916
rect 10068 41914 10092 41916
rect 10148 41914 10154 41916
rect 9908 41862 9910 41914
rect 10090 41862 10092 41914
rect 9846 41860 9852 41862
rect 9908 41860 9932 41862
rect 9988 41860 10012 41862
rect 10068 41860 10092 41862
rect 10148 41860 10154 41862
rect 9846 41840 10154 41860
rect 6880 41372 7188 41392
rect 6880 41370 6886 41372
rect 6942 41370 6966 41372
rect 7022 41370 7046 41372
rect 7102 41370 7126 41372
rect 7182 41370 7188 41372
rect 6942 41318 6944 41370
rect 7124 41318 7126 41370
rect 6880 41316 6886 41318
rect 6942 41316 6966 41318
rect 7022 41316 7046 41318
rect 7102 41316 7126 41318
rect 7182 41316 7188 41318
rect 6880 41296 7188 41316
rect 12811 41372 13119 41392
rect 12811 41370 12817 41372
rect 12873 41370 12897 41372
rect 12953 41370 12977 41372
rect 13033 41370 13057 41372
rect 13113 41370 13119 41372
rect 12873 41318 12875 41370
rect 13055 41318 13057 41370
rect 12811 41316 12817 41318
rect 12873 41316 12897 41318
rect 12953 41316 12977 41318
rect 13033 41316 13057 41318
rect 13113 41316 13119 41318
rect 12811 41296 13119 41316
rect 3915 40828 4223 40848
rect 3915 40826 3921 40828
rect 3977 40826 4001 40828
rect 4057 40826 4081 40828
rect 4137 40826 4161 40828
rect 4217 40826 4223 40828
rect 3977 40774 3979 40826
rect 4159 40774 4161 40826
rect 3915 40772 3921 40774
rect 3977 40772 4001 40774
rect 4057 40772 4081 40774
rect 4137 40772 4161 40774
rect 4217 40772 4223 40774
rect 3915 40752 4223 40772
rect 9846 40828 10154 40848
rect 9846 40826 9852 40828
rect 9908 40826 9932 40828
rect 9988 40826 10012 40828
rect 10068 40826 10092 40828
rect 10148 40826 10154 40828
rect 9908 40774 9910 40826
rect 10090 40774 10092 40826
rect 9846 40772 9852 40774
rect 9908 40772 9932 40774
rect 9988 40772 10012 40774
rect 10068 40772 10092 40774
rect 10148 40772 10154 40774
rect 9846 40752 10154 40772
rect 6880 40284 7188 40304
rect 6880 40282 6886 40284
rect 6942 40282 6966 40284
rect 7022 40282 7046 40284
rect 7102 40282 7126 40284
rect 7182 40282 7188 40284
rect 6942 40230 6944 40282
rect 7124 40230 7126 40282
rect 6880 40228 6886 40230
rect 6942 40228 6966 40230
rect 7022 40228 7046 40230
rect 7102 40228 7126 40230
rect 7182 40228 7188 40230
rect 6880 40208 7188 40228
rect 12811 40284 13119 40304
rect 12811 40282 12817 40284
rect 12873 40282 12897 40284
rect 12953 40282 12977 40284
rect 13033 40282 13057 40284
rect 13113 40282 13119 40284
rect 12873 40230 12875 40282
rect 13055 40230 13057 40282
rect 12811 40228 12817 40230
rect 12873 40228 12897 40230
rect 12953 40228 12977 40230
rect 13033 40228 13057 40230
rect 13113 40228 13119 40230
rect 12811 40208 13119 40228
rect 3915 39740 4223 39760
rect 3915 39738 3921 39740
rect 3977 39738 4001 39740
rect 4057 39738 4081 39740
rect 4137 39738 4161 39740
rect 4217 39738 4223 39740
rect 3977 39686 3979 39738
rect 4159 39686 4161 39738
rect 3915 39684 3921 39686
rect 3977 39684 4001 39686
rect 4057 39684 4081 39686
rect 4137 39684 4161 39686
rect 4217 39684 4223 39686
rect 3915 39664 4223 39684
rect 9846 39740 10154 39760
rect 9846 39738 9852 39740
rect 9908 39738 9932 39740
rect 9988 39738 10012 39740
rect 10068 39738 10092 39740
rect 10148 39738 10154 39740
rect 9908 39686 9910 39738
rect 10090 39686 10092 39738
rect 9846 39684 9852 39686
rect 9908 39684 9932 39686
rect 9988 39684 10012 39686
rect 10068 39684 10092 39686
rect 10148 39684 10154 39686
rect 9846 39664 10154 39684
rect 6880 39196 7188 39216
rect 6880 39194 6886 39196
rect 6942 39194 6966 39196
rect 7022 39194 7046 39196
rect 7102 39194 7126 39196
rect 7182 39194 7188 39196
rect 6942 39142 6944 39194
rect 7124 39142 7126 39194
rect 6880 39140 6886 39142
rect 6942 39140 6966 39142
rect 7022 39140 7046 39142
rect 7102 39140 7126 39142
rect 7182 39140 7188 39142
rect 6880 39120 7188 39140
rect 12811 39196 13119 39216
rect 12811 39194 12817 39196
rect 12873 39194 12897 39196
rect 12953 39194 12977 39196
rect 13033 39194 13057 39196
rect 13113 39194 13119 39196
rect 12873 39142 12875 39194
rect 13055 39142 13057 39194
rect 12811 39140 12817 39142
rect 12873 39140 12897 39142
rect 12953 39140 12977 39142
rect 13033 39140 13057 39142
rect 13113 39140 13119 39142
rect 12811 39120 13119 39140
rect 3915 38652 4223 38672
rect 3915 38650 3921 38652
rect 3977 38650 4001 38652
rect 4057 38650 4081 38652
rect 4137 38650 4161 38652
rect 4217 38650 4223 38652
rect 3977 38598 3979 38650
rect 4159 38598 4161 38650
rect 3915 38596 3921 38598
rect 3977 38596 4001 38598
rect 4057 38596 4081 38598
rect 4137 38596 4161 38598
rect 4217 38596 4223 38598
rect 3915 38576 4223 38596
rect 9846 38652 10154 38672
rect 9846 38650 9852 38652
rect 9908 38650 9932 38652
rect 9988 38650 10012 38652
rect 10068 38650 10092 38652
rect 10148 38650 10154 38652
rect 9908 38598 9910 38650
rect 10090 38598 10092 38650
rect 9846 38596 9852 38598
rect 9908 38596 9932 38598
rect 9988 38596 10012 38598
rect 10068 38596 10092 38598
rect 10148 38596 10154 38598
rect 9846 38576 10154 38596
rect 6880 38108 7188 38128
rect 6880 38106 6886 38108
rect 6942 38106 6966 38108
rect 7022 38106 7046 38108
rect 7102 38106 7126 38108
rect 7182 38106 7188 38108
rect 6942 38054 6944 38106
rect 7124 38054 7126 38106
rect 6880 38052 6886 38054
rect 6942 38052 6966 38054
rect 7022 38052 7046 38054
rect 7102 38052 7126 38054
rect 7182 38052 7188 38054
rect 6880 38032 7188 38052
rect 12811 38108 13119 38128
rect 12811 38106 12817 38108
rect 12873 38106 12897 38108
rect 12953 38106 12977 38108
rect 13033 38106 13057 38108
rect 13113 38106 13119 38108
rect 12873 38054 12875 38106
rect 13055 38054 13057 38106
rect 12811 38052 12817 38054
rect 12873 38052 12897 38054
rect 12953 38052 12977 38054
rect 13033 38052 13057 38054
rect 13113 38052 13119 38054
rect 12811 38032 13119 38052
rect 3915 37564 4223 37584
rect 3915 37562 3921 37564
rect 3977 37562 4001 37564
rect 4057 37562 4081 37564
rect 4137 37562 4161 37564
rect 4217 37562 4223 37564
rect 3977 37510 3979 37562
rect 4159 37510 4161 37562
rect 3915 37508 3921 37510
rect 3977 37508 4001 37510
rect 4057 37508 4081 37510
rect 4137 37508 4161 37510
rect 4217 37508 4223 37510
rect 3915 37488 4223 37508
rect 9846 37564 10154 37584
rect 9846 37562 9852 37564
rect 9908 37562 9932 37564
rect 9988 37562 10012 37564
rect 10068 37562 10092 37564
rect 10148 37562 10154 37564
rect 9908 37510 9910 37562
rect 10090 37510 10092 37562
rect 9846 37508 9852 37510
rect 9908 37508 9932 37510
rect 9988 37508 10012 37510
rect 10068 37508 10092 37510
rect 10148 37508 10154 37510
rect 9846 37488 10154 37508
rect 6880 37020 7188 37040
rect 6880 37018 6886 37020
rect 6942 37018 6966 37020
rect 7022 37018 7046 37020
rect 7102 37018 7126 37020
rect 7182 37018 7188 37020
rect 6942 36966 6944 37018
rect 7124 36966 7126 37018
rect 6880 36964 6886 36966
rect 6942 36964 6966 36966
rect 7022 36964 7046 36966
rect 7102 36964 7126 36966
rect 7182 36964 7188 36966
rect 6880 36944 7188 36964
rect 12811 37020 13119 37040
rect 12811 37018 12817 37020
rect 12873 37018 12897 37020
rect 12953 37018 12977 37020
rect 13033 37018 13057 37020
rect 13113 37018 13119 37020
rect 12873 36966 12875 37018
rect 13055 36966 13057 37018
rect 12811 36964 12817 36966
rect 12873 36964 12897 36966
rect 12953 36964 12977 36966
rect 13033 36964 13057 36966
rect 13113 36964 13119 36966
rect 12811 36944 13119 36964
rect 3915 36476 4223 36496
rect 3915 36474 3921 36476
rect 3977 36474 4001 36476
rect 4057 36474 4081 36476
rect 4137 36474 4161 36476
rect 4217 36474 4223 36476
rect 3977 36422 3979 36474
rect 4159 36422 4161 36474
rect 3915 36420 3921 36422
rect 3977 36420 4001 36422
rect 4057 36420 4081 36422
rect 4137 36420 4161 36422
rect 4217 36420 4223 36422
rect 3915 36400 4223 36420
rect 9846 36476 10154 36496
rect 9846 36474 9852 36476
rect 9908 36474 9932 36476
rect 9988 36474 10012 36476
rect 10068 36474 10092 36476
rect 10148 36474 10154 36476
rect 9908 36422 9910 36474
rect 10090 36422 10092 36474
rect 9846 36420 9852 36422
rect 9908 36420 9932 36422
rect 9988 36420 10012 36422
rect 10068 36420 10092 36422
rect 10148 36420 10154 36422
rect 9846 36400 10154 36420
rect 6880 35932 7188 35952
rect 6880 35930 6886 35932
rect 6942 35930 6966 35932
rect 7022 35930 7046 35932
rect 7102 35930 7126 35932
rect 7182 35930 7188 35932
rect 6942 35878 6944 35930
rect 7124 35878 7126 35930
rect 6880 35876 6886 35878
rect 6942 35876 6966 35878
rect 7022 35876 7046 35878
rect 7102 35876 7126 35878
rect 7182 35876 7188 35878
rect 6880 35856 7188 35876
rect 12811 35932 13119 35952
rect 12811 35930 12817 35932
rect 12873 35930 12897 35932
rect 12953 35930 12977 35932
rect 13033 35930 13057 35932
rect 13113 35930 13119 35932
rect 12873 35878 12875 35930
rect 13055 35878 13057 35930
rect 12811 35876 12817 35878
rect 12873 35876 12897 35878
rect 12953 35876 12977 35878
rect 13033 35876 13057 35878
rect 13113 35876 13119 35878
rect 12811 35856 13119 35876
rect 3915 35388 4223 35408
rect 3915 35386 3921 35388
rect 3977 35386 4001 35388
rect 4057 35386 4081 35388
rect 4137 35386 4161 35388
rect 4217 35386 4223 35388
rect 3977 35334 3979 35386
rect 4159 35334 4161 35386
rect 3915 35332 3921 35334
rect 3977 35332 4001 35334
rect 4057 35332 4081 35334
rect 4137 35332 4161 35334
rect 4217 35332 4223 35334
rect 3915 35312 4223 35332
rect 9846 35388 10154 35408
rect 9846 35386 9852 35388
rect 9908 35386 9932 35388
rect 9988 35386 10012 35388
rect 10068 35386 10092 35388
rect 10148 35386 10154 35388
rect 9908 35334 9910 35386
rect 10090 35334 10092 35386
rect 9846 35332 9852 35334
rect 9908 35332 9932 35334
rect 9988 35332 10012 35334
rect 10068 35332 10092 35334
rect 10148 35332 10154 35334
rect 9846 35312 10154 35332
rect 2044 35012 2096 35018
rect 2044 34954 2096 34960
rect 6880 34844 7188 34864
rect 6880 34842 6886 34844
rect 6942 34842 6966 34844
rect 7022 34842 7046 34844
rect 7102 34842 7126 34844
rect 7182 34842 7188 34844
rect 6942 34790 6944 34842
rect 7124 34790 7126 34842
rect 6880 34788 6886 34790
rect 6942 34788 6966 34790
rect 7022 34788 7046 34790
rect 7102 34788 7126 34790
rect 7182 34788 7188 34790
rect 6880 34768 7188 34788
rect 12811 34844 13119 34864
rect 12811 34842 12817 34844
rect 12873 34842 12897 34844
rect 12953 34842 12977 34844
rect 13033 34842 13057 34844
rect 13113 34842 13119 34844
rect 12873 34790 12875 34842
rect 13055 34790 13057 34842
rect 12811 34788 12817 34790
rect 12873 34788 12897 34790
rect 12953 34788 12977 34790
rect 13033 34788 13057 34790
rect 13113 34788 13119 34790
rect 12811 34768 13119 34788
rect 13636 34468 13688 34474
rect 13636 34410 13688 34416
rect 13452 34400 13504 34406
rect 13452 34342 13504 34348
rect 3915 34300 4223 34320
rect 3915 34298 3921 34300
rect 3977 34298 4001 34300
rect 4057 34298 4081 34300
rect 4137 34298 4161 34300
rect 4217 34298 4223 34300
rect 3977 34246 3979 34298
rect 4159 34246 4161 34298
rect 3915 34244 3921 34246
rect 3977 34244 4001 34246
rect 4057 34244 4081 34246
rect 4137 34244 4161 34246
rect 4217 34244 4223 34246
rect 3915 34224 4223 34244
rect 9846 34300 10154 34320
rect 9846 34298 9852 34300
rect 9908 34298 9932 34300
rect 9988 34298 10012 34300
rect 10068 34298 10092 34300
rect 10148 34298 10154 34300
rect 9908 34246 9910 34298
rect 10090 34246 10092 34298
rect 9846 34244 9852 34246
rect 9908 34244 9932 34246
rect 9988 34244 10012 34246
rect 10068 34244 10092 34246
rect 10148 34244 10154 34246
rect 9846 34224 10154 34244
rect 13464 34202 13492 34342
rect 13452 34196 13504 34202
rect 13452 34138 13504 34144
rect 13648 34066 13676 34410
rect 13636 34060 13688 34066
rect 13636 34002 13688 34008
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 13452 33856 13504 33862
rect 13452 33798 13504 33804
rect 6880 33756 7188 33776
rect 6880 33754 6886 33756
rect 6942 33754 6966 33756
rect 7022 33754 7046 33756
rect 7102 33754 7126 33756
rect 7182 33754 7188 33756
rect 6942 33702 6944 33754
rect 7124 33702 7126 33754
rect 6880 33700 6886 33702
rect 6942 33700 6966 33702
rect 7022 33700 7046 33702
rect 7102 33700 7126 33702
rect 7182 33700 7188 33702
rect 6880 33680 7188 33700
rect 3915 33212 4223 33232
rect 3915 33210 3921 33212
rect 3977 33210 4001 33212
rect 4057 33210 4081 33212
rect 4137 33210 4161 33212
rect 4217 33210 4223 33212
rect 3977 33158 3979 33210
rect 4159 33158 4161 33210
rect 3915 33156 3921 33158
rect 3977 33156 4001 33158
rect 4057 33156 4081 33158
rect 4137 33156 4161 33158
rect 4217 33156 4223 33158
rect 3915 33136 4223 33156
rect 9846 33212 10154 33232
rect 9846 33210 9852 33212
rect 9908 33210 9932 33212
rect 9988 33210 10012 33212
rect 10068 33210 10092 33212
rect 10148 33210 10154 33212
rect 9908 33158 9910 33210
rect 10090 33158 10092 33210
rect 9846 33156 9852 33158
rect 9908 33156 9932 33158
rect 9988 33156 10012 33158
rect 10068 33156 10092 33158
rect 10148 33156 10154 33158
rect 9846 33136 10154 33156
rect 12728 32774 12756 33798
rect 12811 33756 13119 33776
rect 12811 33754 12817 33756
rect 12873 33754 12897 33756
rect 12953 33754 12977 33756
rect 13033 33754 13057 33756
rect 13113 33754 13119 33756
rect 12873 33702 12875 33754
rect 13055 33702 13057 33754
rect 12811 33700 12817 33702
rect 12873 33700 12897 33702
rect 12953 33700 12977 33702
rect 13033 33700 13057 33702
rect 13113 33700 13119 33702
rect 12811 33680 13119 33700
rect 13464 33522 13492 33798
rect 13542 33552 13598 33561
rect 13452 33516 13504 33522
rect 13542 33487 13544 33496
rect 13452 33458 13504 33464
rect 13596 33487 13598 33496
rect 13544 33458 13596 33464
rect 12716 32768 12768 32774
rect 12716 32710 12768 32716
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 6880 32668 7188 32688
rect 6880 32666 6886 32668
rect 6942 32666 6966 32668
rect 7022 32666 7046 32668
rect 7102 32666 7126 32668
rect 7182 32666 7188 32668
rect 6942 32614 6944 32666
rect 7124 32614 7126 32666
rect 6880 32612 6886 32614
rect 6942 32612 6966 32614
rect 7022 32612 7046 32614
rect 7102 32612 7126 32614
rect 7182 32612 7188 32614
rect 6880 32592 7188 32612
rect 3915 32124 4223 32144
rect 3915 32122 3921 32124
rect 3977 32122 4001 32124
rect 4057 32122 4081 32124
rect 4137 32122 4161 32124
rect 4217 32122 4223 32124
rect 3977 32070 3979 32122
rect 4159 32070 4161 32122
rect 3915 32068 3921 32070
rect 3977 32068 4001 32070
rect 4057 32068 4081 32070
rect 4137 32068 4161 32070
rect 4217 32068 4223 32070
rect 3915 32048 4223 32068
rect 9846 32124 10154 32144
rect 9846 32122 9852 32124
rect 9908 32122 9932 32124
rect 9988 32122 10012 32124
rect 10068 32122 10092 32124
rect 10148 32122 10154 32124
rect 9908 32070 9910 32122
rect 10090 32070 10092 32122
rect 9846 32068 9852 32070
rect 9908 32068 9932 32070
rect 9988 32068 10012 32070
rect 10068 32068 10092 32070
rect 10148 32068 10154 32070
rect 9846 32048 10154 32068
rect 6880 31580 7188 31600
rect 6880 31578 6886 31580
rect 6942 31578 6966 31580
rect 7022 31578 7046 31580
rect 7102 31578 7126 31580
rect 7182 31578 7188 31580
rect 6942 31526 6944 31578
rect 7124 31526 7126 31578
rect 6880 31524 6886 31526
rect 6942 31524 6966 31526
rect 7022 31524 7046 31526
rect 7102 31524 7126 31526
rect 7182 31524 7188 31526
rect 6880 31504 7188 31524
rect 12728 31414 12756 32710
rect 12811 32668 13119 32688
rect 12811 32666 12817 32668
rect 12873 32666 12897 32668
rect 12953 32666 12977 32668
rect 13033 32666 13057 32668
rect 13113 32666 13119 32668
rect 12873 32614 12875 32666
rect 13055 32614 13057 32666
rect 12811 32612 12817 32614
rect 12873 32612 12897 32614
rect 12953 32612 12977 32614
rect 13033 32612 13057 32614
rect 13113 32612 13119 32614
rect 12811 32592 13119 32612
rect 13372 31822 13400 32710
rect 13648 32570 13676 34002
rect 13636 32564 13688 32570
rect 13636 32506 13688 32512
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 12811 31580 13119 31600
rect 12811 31578 12817 31580
rect 12873 31578 12897 31580
rect 12953 31578 12977 31580
rect 13033 31578 13057 31580
rect 13113 31578 13119 31580
rect 12873 31526 12875 31578
rect 13055 31526 13057 31578
rect 12811 31524 12817 31526
rect 12873 31524 12897 31526
rect 12953 31524 12977 31526
rect 13033 31524 13057 31526
rect 13113 31524 13119 31526
rect 12811 31504 13119 31524
rect 12716 31408 12768 31414
rect 12716 31350 12768 31356
rect 3915 31036 4223 31056
rect 3915 31034 3921 31036
rect 3977 31034 4001 31036
rect 4057 31034 4081 31036
rect 4137 31034 4161 31036
rect 4217 31034 4223 31036
rect 3977 30982 3979 31034
rect 4159 30982 4161 31034
rect 3915 30980 3921 30982
rect 3977 30980 4001 30982
rect 4057 30980 4081 30982
rect 4137 30980 4161 30982
rect 4217 30980 4223 30982
rect 3915 30960 4223 30980
rect 9846 31036 10154 31056
rect 9846 31034 9852 31036
rect 9908 31034 9932 31036
rect 9988 31034 10012 31036
rect 10068 31034 10092 31036
rect 10148 31034 10154 31036
rect 9908 30982 9910 31034
rect 10090 30982 10092 31034
rect 9846 30980 9852 30982
rect 9908 30980 9932 30982
rect 9988 30980 10012 30982
rect 10068 30980 10092 30982
rect 10148 30980 10154 30982
rect 9846 30960 10154 30980
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 30569 1440 30670
rect 1398 30560 1454 30569
rect 1398 30495 1454 30504
rect 1412 30394 1440 30495
rect 6880 30492 7188 30512
rect 6880 30490 6886 30492
rect 6942 30490 6966 30492
rect 7022 30490 7046 30492
rect 7102 30490 7126 30492
rect 7182 30490 7188 30492
rect 6942 30438 6944 30490
rect 7124 30438 7126 30490
rect 6880 30436 6886 30438
rect 6942 30436 6966 30438
rect 7022 30436 7046 30438
rect 7102 30436 7126 30438
rect 7182 30436 7188 30438
rect 6880 30416 7188 30436
rect 1400 30388 1452 30394
rect 1400 30330 1452 30336
rect 3915 29948 4223 29968
rect 3915 29946 3921 29948
rect 3977 29946 4001 29948
rect 4057 29946 4081 29948
rect 4137 29946 4161 29948
rect 4217 29946 4223 29948
rect 3977 29894 3979 29946
rect 4159 29894 4161 29946
rect 3915 29892 3921 29894
rect 3977 29892 4001 29894
rect 4057 29892 4081 29894
rect 4137 29892 4161 29894
rect 4217 29892 4223 29894
rect 3915 29872 4223 29892
rect 9846 29948 10154 29968
rect 9846 29946 9852 29948
rect 9908 29946 9932 29948
rect 9988 29946 10012 29948
rect 10068 29946 10092 29948
rect 10148 29946 10154 29948
rect 9908 29894 9910 29946
rect 10090 29894 10092 29946
rect 9846 29892 9852 29894
rect 9908 29892 9932 29894
rect 9988 29892 10012 29894
rect 10068 29892 10092 29894
rect 10148 29892 10154 29894
rect 9846 29872 10154 29892
rect 6880 29404 7188 29424
rect 6880 29402 6886 29404
rect 6942 29402 6966 29404
rect 7022 29402 7046 29404
rect 7102 29402 7126 29404
rect 7182 29402 7188 29404
rect 6942 29350 6944 29402
rect 7124 29350 7126 29402
rect 6880 29348 6886 29350
rect 6942 29348 6966 29350
rect 7022 29348 7046 29350
rect 7102 29348 7126 29350
rect 7182 29348 7188 29350
rect 6880 29328 7188 29348
rect 3915 28860 4223 28880
rect 3915 28858 3921 28860
rect 3977 28858 4001 28860
rect 4057 28858 4081 28860
rect 4137 28858 4161 28860
rect 4217 28858 4223 28860
rect 3977 28806 3979 28858
rect 4159 28806 4161 28858
rect 3915 28804 3921 28806
rect 3977 28804 4001 28806
rect 4057 28804 4081 28806
rect 4137 28804 4161 28806
rect 4217 28804 4223 28806
rect 3915 28784 4223 28804
rect 9846 28860 10154 28880
rect 9846 28858 9852 28860
rect 9908 28858 9932 28860
rect 9988 28858 10012 28860
rect 10068 28858 10092 28860
rect 10148 28858 10154 28860
rect 9908 28806 9910 28858
rect 10090 28806 10092 28858
rect 9846 28804 9852 28806
rect 9908 28804 9932 28806
rect 9988 28804 10012 28806
rect 10068 28804 10092 28806
rect 10148 28804 10154 28806
rect 9846 28784 10154 28804
rect 6880 28316 7188 28336
rect 6880 28314 6886 28316
rect 6942 28314 6966 28316
rect 7022 28314 7046 28316
rect 7102 28314 7126 28316
rect 7182 28314 7188 28316
rect 6942 28262 6944 28314
rect 7124 28262 7126 28314
rect 6880 28260 6886 28262
rect 6942 28260 6966 28262
rect 7022 28260 7046 28262
rect 7102 28260 7126 28262
rect 7182 28260 7188 28262
rect 6880 28240 7188 28260
rect 3915 27772 4223 27792
rect 3915 27770 3921 27772
rect 3977 27770 4001 27772
rect 4057 27770 4081 27772
rect 4137 27770 4161 27772
rect 4217 27770 4223 27772
rect 3977 27718 3979 27770
rect 4159 27718 4161 27770
rect 3915 27716 3921 27718
rect 3977 27716 4001 27718
rect 4057 27716 4081 27718
rect 4137 27716 4161 27718
rect 4217 27716 4223 27718
rect 3915 27696 4223 27716
rect 9846 27772 10154 27792
rect 9846 27770 9852 27772
rect 9908 27770 9932 27772
rect 9988 27770 10012 27772
rect 10068 27770 10092 27772
rect 10148 27770 10154 27772
rect 9908 27718 9910 27770
rect 10090 27718 10092 27770
rect 9846 27716 9852 27718
rect 9908 27716 9932 27718
rect 9988 27716 10012 27718
rect 10068 27716 10092 27718
rect 10148 27716 10154 27718
rect 9846 27696 10154 27716
rect 6880 27228 7188 27248
rect 6880 27226 6886 27228
rect 6942 27226 6966 27228
rect 7022 27226 7046 27228
rect 7102 27226 7126 27228
rect 7182 27226 7188 27228
rect 6942 27174 6944 27226
rect 7124 27174 7126 27226
rect 6880 27172 6886 27174
rect 6942 27172 6966 27174
rect 7022 27172 7046 27174
rect 7102 27172 7126 27174
rect 7182 27172 7188 27174
rect 6880 27152 7188 27172
rect 3915 26684 4223 26704
rect 3915 26682 3921 26684
rect 3977 26682 4001 26684
rect 4057 26682 4081 26684
rect 4137 26682 4161 26684
rect 4217 26682 4223 26684
rect 3977 26630 3979 26682
rect 4159 26630 4161 26682
rect 3915 26628 3921 26630
rect 3977 26628 4001 26630
rect 4057 26628 4081 26630
rect 4137 26628 4161 26630
rect 4217 26628 4223 26630
rect 3915 26608 4223 26628
rect 9846 26684 10154 26704
rect 9846 26682 9852 26684
rect 9908 26682 9932 26684
rect 9988 26682 10012 26684
rect 10068 26682 10092 26684
rect 10148 26682 10154 26684
rect 9908 26630 9910 26682
rect 10090 26630 10092 26682
rect 9846 26628 9852 26630
rect 9908 26628 9932 26630
rect 9988 26628 10012 26630
rect 10068 26628 10092 26630
rect 10148 26628 10154 26630
rect 9846 26608 10154 26628
rect 6880 26140 7188 26160
rect 6880 26138 6886 26140
rect 6942 26138 6966 26140
rect 7022 26138 7046 26140
rect 7102 26138 7126 26140
rect 7182 26138 7188 26140
rect 6942 26086 6944 26138
rect 7124 26086 7126 26138
rect 6880 26084 6886 26086
rect 6942 26084 6966 26086
rect 7022 26084 7046 26086
rect 7102 26084 7126 26086
rect 7182 26084 7188 26086
rect 6880 26064 7188 26084
rect 3915 25596 4223 25616
rect 3915 25594 3921 25596
rect 3977 25594 4001 25596
rect 4057 25594 4081 25596
rect 4137 25594 4161 25596
rect 4217 25594 4223 25596
rect 3977 25542 3979 25594
rect 4159 25542 4161 25594
rect 3915 25540 3921 25542
rect 3977 25540 4001 25542
rect 4057 25540 4081 25542
rect 4137 25540 4161 25542
rect 4217 25540 4223 25542
rect 3915 25520 4223 25540
rect 9846 25596 10154 25616
rect 9846 25594 9852 25596
rect 9908 25594 9932 25596
rect 9988 25594 10012 25596
rect 10068 25594 10092 25596
rect 10148 25594 10154 25596
rect 9908 25542 9910 25594
rect 10090 25542 10092 25594
rect 9846 25540 9852 25542
rect 9908 25540 9932 25542
rect 9988 25540 10012 25542
rect 10068 25540 10092 25542
rect 10148 25540 10154 25542
rect 9846 25520 10154 25540
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1504 24993 1532 25094
rect 6880 25052 7188 25072
rect 6880 25050 6886 25052
rect 6942 25050 6966 25052
rect 7022 25050 7046 25052
rect 7102 25050 7126 25052
rect 7182 25050 7188 25052
rect 6942 24998 6944 25050
rect 7124 24998 7126 25050
rect 6880 24996 6886 24998
rect 6942 24996 6966 24998
rect 7022 24996 7046 24998
rect 7102 24996 7126 24998
rect 7182 24996 7188 24998
rect 1490 24984 1546 24993
rect 6880 24976 7188 24996
rect 1490 24919 1546 24928
rect 1676 24812 1728 24818
rect 1676 24754 1728 24760
rect 1688 19922 1716 24754
rect 3915 24508 4223 24528
rect 3915 24506 3921 24508
rect 3977 24506 4001 24508
rect 4057 24506 4081 24508
rect 4137 24506 4161 24508
rect 4217 24506 4223 24508
rect 3977 24454 3979 24506
rect 4159 24454 4161 24506
rect 3915 24452 3921 24454
rect 3977 24452 4001 24454
rect 4057 24452 4081 24454
rect 4137 24452 4161 24454
rect 4217 24452 4223 24454
rect 3915 24432 4223 24452
rect 9846 24508 10154 24528
rect 9846 24506 9852 24508
rect 9908 24506 9932 24508
rect 9988 24506 10012 24508
rect 10068 24506 10092 24508
rect 10148 24506 10154 24508
rect 9908 24454 9910 24506
rect 10090 24454 10092 24506
rect 9846 24452 9852 24454
rect 9908 24452 9932 24454
rect 9988 24452 10012 24454
rect 10068 24452 10092 24454
rect 10148 24452 10154 24454
rect 9846 24432 10154 24452
rect 11164 24342 11192 25230
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 11152 24336 11204 24342
rect 11152 24278 11204 24284
rect 12544 24206 12572 24754
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 6880 23964 7188 23984
rect 6880 23962 6886 23964
rect 6942 23962 6966 23964
rect 7022 23962 7046 23964
rect 7102 23962 7126 23964
rect 7182 23962 7188 23964
rect 6942 23910 6944 23962
rect 7124 23910 7126 23962
rect 6880 23908 6886 23910
rect 6942 23908 6966 23910
rect 7022 23908 7046 23910
rect 7102 23908 7126 23910
rect 7182 23908 7188 23910
rect 6880 23888 7188 23908
rect 3915 23420 4223 23440
rect 3915 23418 3921 23420
rect 3977 23418 4001 23420
rect 4057 23418 4081 23420
rect 4137 23418 4161 23420
rect 4217 23418 4223 23420
rect 3977 23366 3979 23418
rect 4159 23366 4161 23418
rect 3915 23364 3921 23366
rect 3977 23364 4001 23366
rect 4057 23364 4081 23366
rect 4137 23364 4161 23366
rect 4217 23364 4223 23366
rect 3915 23344 4223 23364
rect 9846 23420 10154 23440
rect 9846 23418 9852 23420
rect 9908 23418 9932 23420
rect 9988 23418 10012 23420
rect 10068 23418 10092 23420
rect 10148 23418 10154 23420
rect 9908 23366 9910 23418
rect 10090 23366 10092 23418
rect 9846 23364 9852 23366
rect 9908 23364 9932 23366
rect 9988 23364 10012 23366
rect 10068 23364 10092 23366
rect 10148 23364 10154 23366
rect 9846 23344 10154 23364
rect 6880 22876 7188 22896
rect 6880 22874 6886 22876
rect 6942 22874 6966 22876
rect 7022 22874 7046 22876
rect 7102 22874 7126 22876
rect 7182 22874 7188 22876
rect 6942 22822 6944 22874
rect 7124 22822 7126 22874
rect 6880 22820 6886 22822
rect 6942 22820 6966 22822
rect 7022 22820 7046 22822
rect 7102 22820 7126 22822
rect 7182 22820 7188 22822
rect 6880 22800 7188 22820
rect 3915 22332 4223 22352
rect 3915 22330 3921 22332
rect 3977 22330 4001 22332
rect 4057 22330 4081 22332
rect 4137 22330 4161 22332
rect 4217 22330 4223 22332
rect 3977 22278 3979 22330
rect 4159 22278 4161 22330
rect 3915 22276 3921 22278
rect 3977 22276 4001 22278
rect 4057 22276 4081 22278
rect 4137 22276 4161 22278
rect 4217 22276 4223 22278
rect 3915 22256 4223 22276
rect 9846 22332 10154 22352
rect 9846 22330 9852 22332
rect 9908 22330 9932 22332
rect 9988 22330 10012 22332
rect 10068 22330 10092 22332
rect 10148 22330 10154 22332
rect 9908 22278 9910 22330
rect 10090 22278 10092 22330
rect 9846 22276 9852 22278
rect 9908 22276 9932 22278
rect 9988 22276 10012 22278
rect 10068 22276 10092 22278
rect 10148 22276 10154 22278
rect 9846 22256 10154 22276
rect 6880 21788 7188 21808
rect 6880 21786 6886 21788
rect 6942 21786 6966 21788
rect 7022 21786 7046 21788
rect 7102 21786 7126 21788
rect 7182 21786 7188 21788
rect 6942 21734 6944 21786
rect 7124 21734 7126 21786
rect 6880 21732 6886 21734
rect 6942 21732 6966 21734
rect 7022 21732 7046 21734
rect 7102 21732 7126 21734
rect 7182 21732 7188 21734
rect 6880 21712 7188 21732
rect 3915 21244 4223 21264
rect 3915 21242 3921 21244
rect 3977 21242 4001 21244
rect 4057 21242 4081 21244
rect 4137 21242 4161 21244
rect 4217 21242 4223 21244
rect 3977 21190 3979 21242
rect 4159 21190 4161 21242
rect 3915 21188 3921 21190
rect 3977 21188 4001 21190
rect 4057 21188 4081 21190
rect 4137 21188 4161 21190
rect 4217 21188 4223 21190
rect 3915 21168 4223 21188
rect 9846 21244 10154 21264
rect 9846 21242 9852 21244
rect 9908 21242 9932 21244
rect 9988 21242 10012 21244
rect 10068 21242 10092 21244
rect 10148 21242 10154 21244
rect 9908 21190 9910 21242
rect 10090 21190 10092 21242
rect 9846 21188 9852 21190
rect 9908 21188 9932 21190
rect 9988 21188 10012 21190
rect 10068 21188 10092 21190
rect 10148 21188 10154 21190
rect 9846 21168 10154 21188
rect 6880 20700 7188 20720
rect 6880 20698 6886 20700
rect 6942 20698 6966 20700
rect 7022 20698 7046 20700
rect 7102 20698 7126 20700
rect 7182 20698 7188 20700
rect 6942 20646 6944 20698
rect 7124 20646 7126 20698
rect 6880 20644 6886 20646
rect 6942 20644 6966 20646
rect 7022 20644 7046 20646
rect 7102 20644 7126 20646
rect 7182 20644 7188 20646
rect 6880 20624 7188 20644
rect 3915 20156 4223 20176
rect 3915 20154 3921 20156
rect 3977 20154 4001 20156
rect 4057 20154 4081 20156
rect 4137 20154 4161 20156
rect 4217 20154 4223 20156
rect 3977 20102 3979 20154
rect 4159 20102 4161 20154
rect 3915 20100 3921 20102
rect 3977 20100 4001 20102
rect 4057 20100 4081 20102
rect 4137 20100 4161 20102
rect 4217 20100 4223 20102
rect 3915 20080 4223 20100
rect 9846 20156 10154 20176
rect 9846 20154 9852 20156
rect 9908 20154 9932 20156
rect 9988 20154 10012 20156
rect 10068 20154 10092 20156
rect 10148 20154 10154 20156
rect 9908 20102 9910 20154
rect 10090 20102 10092 20154
rect 9846 20100 9852 20102
rect 9908 20100 9932 20102
rect 9988 20100 10012 20102
rect 10068 20100 10092 20102
rect 10148 20100 10154 20102
rect 9846 20080 10154 20100
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1412 19446 1440 19790
rect 6880 19612 7188 19632
rect 6880 19610 6886 19612
rect 6942 19610 6966 19612
rect 7022 19610 7046 19612
rect 7102 19610 7126 19612
rect 7182 19610 7188 19612
rect 6942 19558 6944 19610
rect 7124 19558 7126 19610
rect 6880 19556 6886 19558
rect 6942 19556 6966 19558
rect 7022 19556 7046 19558
rect 7102 19556 7126 19558
rect 7182 19556 7188 19558
rect 6880 19536 7188 19556
rect 1400 19440 1452 19446
rect 1398 19408 1400 19417
rect 1452 19408 1454 19417
rect 1398 19343 1454 19352
rect 3915 19068 4223 19088
rect 3915 19066 3921 19068
rect 3977 19066 4001 19068
rect 4057 19066 4081 19068
rect 4137 19066 4161 19068
rect 4217 19066 4223 19068
rect 3977 19014 3979 19066
rect 4159 19014 4161 19066
rect 3915 19012 3921 19014
rect 3977 19012 4001 19014
rect 4057 19012 4081 19014
rect 4137 19012 4161 19014
rect 4217 19012 4223 19014
rect 3915 18992 4223 19012
rect 9846 19068 10154 19088
rect 9846 19066 9852 19068
rect 9908 19066 9932 19068
rect 9988 19066 10012 19068
rect 10068 19066 10092 19068
rect 10148 19066 10154 19068
rect 9908 19014 9910 19066
rect 10090 19014 10092 19066
rect 9846 19012 9852 19014
rect 9908 19012 9932 19014
rect 9988 19012 10012 19014
rect 10068 19012 10092 19014
rect 10148 19012 10154 19014
rect 9846 18992 10154 19012
rect 6880 18524 7188 18544
rect 6880 18522 6886 18524
rect 6942 18522 6966 18524
rect 7022 18522 7046 18524
rect 7102 18522 7126 18524
rect 7182 18522 7188 18524
rect 6942 18470 6944 18522
rect 7124 18470 7126 18522
rect 6880 18468 6886 18470
rect 6942 18468 6966 18470
rect 7022 18468 7046 18470
rect 7102 18468 7126 18470
rect 7182 18468 7188 18470
rect 6880 18448 7188 18468
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 3915 17980 4223 18000
rect 3915 17978 3921 17980
rect 3977 17978 4001 17980
rect 4057 17978 4081 17980
rect 4137 17978 4161 17980
rect 4217 17978 4223 17980
rect 3977 17926 3979 17978
rect 4159 17926 4161 17978
rect 3915 17924 3921 17926
rect 3977 17924 4001 17926
rect 4057 17924 4081 17926
rect 4137 17924 4161 17926
rect 4217 17924 4223 17926
rect 3915 17904 4223 17924
rect 6880 17436 7188 17456
rect 6880 17434 6886 17436
rect 6942 17434 6966 17436
rect 7022 17434 7046 17436
rect 7102 17434 7126 17436
rect 7182 17434 7188 17436
rect 6942 17382 6944 17434
rect 7124 17382 7126 17434
rect 6880 17380 6886 17382
rect 6942 17380 6966 17382
rect 7022 17380 7046 17382
rect 7102 17380 7126 17382
rect 7182 17380 7188 17382
rect 6880 17360 7188 17380
rect 3915 16892 4223 16912
rect 3915 16890 3921 16892
rect 3977 16890 4001 16892
rect 4057 16890 4081 16892
rect 4137 16890 4161 16892
rect 4217 16890 4223 16892
rect 3977 16838 3979 16890
rect 4159 16838 4161 16890
rect 3915 16836 3921 16838
rect 3977 16836 4001 16838
rect 4057 16836 4081 16838
rect 4137 16836 4161 16838
rect 4217 16836 4223 16838
rect 3915 16816 4223 16836
rect 6880 16348 7188 16368
rect 6880 16346 6886 16348
rect 6942 16346 6966 16348
rect 7022 16346 7046 16348
rect 7102 16346 7126 16348
rect 7182 16346 7188 16348
rect 6942 16294 6944 16346
rect 7124 16294 7126 16346
rect 6880 16292 6886 16294
rect 6942 16292 6966 16294
rect 7022 16292 7046 16294
rect 7102 16292 7126 16294
rect 7182 16292 7188 16294
rect 6880 16272 7188 16292
rect 3915 15804 4223 15824
rect 3915 15802 3921 15804
rect 3977 15802 4001 15804
rect 4057 15802 4081 15804
rect 4137 15802 4161 15804
rect 4217 15802 4223 15804
rect 3977 15750 3979 15802
rect 4159 15750 4161 15802
rect 3915 15748 3921 15750
rect 3977 15748 4001 15750
rect 4057 15748 4081 15750
rect 4137 15748 4161 15750
rect 4217 15748 4223 15750
rect 3915 15728 4223 15748
rect 6880 15260 7188 15280
rect 6880 15258 6886 15260
rect 6942 15258 6966 15260
rect 7022 15258 7046 15260
rect 7102 15258 7126 15260
rect 7182 15258 7188 15260
rect 6942 15206 6944 15258
rect 7124 15206 7126 15258
rect 6880 15204 6886 15206
rect 6942 15204 6966 15206
rect 7022 15204 7046 15206
rect 7102 15204 7126 15206
rect 7182 15204 7188 15206
rect 6880 15184 7188 15204
rect 3915 14716 4223 14736
rect 3915 14714 3921 14716
rect 3977 14714 4001 14716
rect 4057 14714 4081 14716
rect 4137 14714 4161 14716
rect 4217 14714 4223 14716
rect 3977 14662 3979 14714
rect 4159 14662 4161 14714
rect 3915 14660 3921 14662
rect 3977 14660 4001 14662
rect 4057 14660 4081 14662
rect 4137 14660 4161 14662
rect 4217 14660 4223 14662
rect 3915 14640 4223 14660
rect 6880 14172 7188 14192
rect 6880 14170 6886 14172
rect 6942 14170 6966 14172
rect 7022 14170 7046 14172
rect 7102 14170 7126 14172
rect 7182 14170 7188 14172
rect 6942 14118 6944 14170
rect 7124 14118 7126 14170
rect 6880 14116 6886 14118
rect 6942 14116 6966 14118
rect 7022 14116 7046 14118
rect 7102 14116 7126 14118
rect 7182 14116 7188 14118
rect 6880 14096 7188 14116
rect 8312 13938 8340 18158
rect 9846 17980 10154 18000
rect 9846 17978 9852 17980
rect 9908 17978 9932 17980
rect 9988 17978 10012 17980
rect 10068 17978 10092 17980
rect 10148 17978 10154 17980
rect 9908 17926 9910 17978
rect 10090 17926 10092 17978
rect 9846 17924 9852 17926
rect 9908 17924 9932 17926
rect 9988 17924 10012 17926
rect 10068 17924 10092 17926
rect 10148 17924 10154 17926
rect 9846 17904 10154 17924
rect 11348 17542 11376 18226
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 9846 16892 10154 16912
rect 9846 16890 9852 16892
rect 9908 16890 9932 16892
rect 9988 16890 10012 16892
rect 10068 16890 10092 16892
rect 10148 16890 10154 16892
rect 9908 16838 9910 16890
rect 10090 16838 10092 16890
rect 9846 16836 9852 16838
rect 9908 16836 9932 16838
rect 9988 16836 10012 16838
rect 10068 16836 10092 16838
rect 10148 16836 10154 16838
rect 9846 16816 10154 16836
rect 9846 15804 10154 15824
rect 9846 15802 9852 15804
rect 9908 15802 9932 15804
rect 9988 15802 10012 15804
rect 10068 15802 10092 15804
rect 10148 15802 10154 15804
rect 9908 15750 9910 15802
rect 10090 15750 10092 15802
rect 9846 15748 9852 15750
rect 9908 15748 9932 15750
rect 9988 15748 10012 15750
rect 10068 15748 10092 15750
rect 10148 15748 10154 15750
rect 9846 15728 10154 15748
rect 9846 14716 10154 14736
rect 9846 14714 9852 14716
rect 9908 14714 9932 14716
rect 9988 14714 10012 14716
rect 10068 14714 10092 14716
rect 10148 14714 10154 14716
rect 9908 14662 9910 14714
rect 10090 14662 10092 14714
rect 9846 14660 9852 14662
rect 9908 14660 9932 14662
rect 9988 14660 10012 14662
rect 10068 14660 10092 14662
rect 10148 14660 10154 14662
rect 9846 14640 10154 14660
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 1400 13864 1452 13870
rect 1398 13832 1400 13841
rect 1452 13832 1454 13841
rect 1398 13767 1454 13776
rect 1412 13530 1440 13767
rect 3915 13628 4223 13648
rect 3915 13626 3921 13628
rect 3977 13626 4001 13628
rect 4057 13626 4081 13628
rect 4137 13626 4161 13628
rect 4217 13626 4223 13628
rect 3977 13574 3979 13626
rect 4159 13574 4161 13626
rect 3915 13572 3921 13574
rect 3977 13572 4001 13574
rect 4057 13572 4081 13574
rect 4137 13572 4161 13574
rect 4217 13572 4223 13574
rect 3915 13552 4223 13572
rect 9846 13628 10154 13648
rect 9846 13626 9852 13628
rect 9908 13626 9932 13628
rect 9988 13626 10012 13628
rect 10068 13626 10092 13628
rect 10148 13626 10154 13628
rect 9908 13574 9910 13626
rect 10090 13574 10092 13626
rect 9846 13572 9852 13574
rect 9908 13572 9932 13574
rect 9988 13572 10012 13574
rect 10068 13572 10092 13574
rect 10148 13572 10154 13574
rect 9846 13552 10154 13572
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 6880 13084 7188 13104
rect 6880 13082 6886 13084
rect 6942 13082 6966 13084
rect 7022 13082 7046 13084
rect 7102 13082 7126 13084
rect 7182 13082 7188 13084
rect 6942 13030 6944 13082
rect 7124 13030 7126 13082
rect 6880 13028 6886 13030
rect 6942 13028 6966 13030
rect 7022 13028 7046 13030
rect 7102 13028 7126 13030
rect 7182 13028 7188 13030
rect 6880 13008 7188 13028
rect 3915 12540 4223 12560
rect 3915 12538 3921 12540
rect 3977 12538 4001 12540
rect 4057 12538 4081 12540
rect 4137 12538 4161 12540
rect 4217 12538 4223 12540
rect 3977 12486 3979 12538
rect 4159 12486 4161 12538
rect 3915 12484 3921 12486
rect 3977 12484 4001 12486
rect 4057 12484 4081 12486
rect 4137 12484 4161 12486
rect 4217 12484 4223 12486
rect 3915 12464 4223 12484
rect 9846 12540 10154 12560
rect 9846 12538 9852 12540
rect 9908 12538 9932 12540
rect 9988 12538 10012 12540
rect 10068 12538 10092 12540
rect 10148 12538 10154 12540
rect 9908 12486 9910 12538
rect 10090 12486 10092 12538
rect 9846 12484 9852 12486
rect 9908 12484 9932 12486
rect 9988 12484 10012 12486
rect 10068 12484 10092 12486
rect 10148 12484 10154 12486
rect 9846 12464 10154 12484
rect 6880 11996 7188 12016
rect 6880 11994 6886 11996
rect 6942 11994 6966 11996
rect 7022 11994 7046 11996
rect 7102 11994 7126 11996
rect 7182 11994 7188 11996
rect 6942 11942 6944 11994
rect 7124 11942 7126 11994
rect 6880 11940 6886 11942
rect 6942 11940 6966 11942
rect 7022 11940 7046 11942
rect 7102 11940 7126 11942
rect 7182 11940 7188 11942
rect 6880 11920 7188 11940
rect 3915 11452 4223 11472
rect 3915 11450 3921 11452
rect 3977 11450 4001 11452
rect 4057 11450 4081 11452
rect 4137 11450 4161 11452
rect 4217 11450 4223 11452
rect 3977 11398 3979 11450
rect 4159 11398 4161 11450
rect 3915 11396 3921 11398
rect 3977 11396 4001 11398
rect 4057 11396 4081 11398
rect 4137 11396 4161 11398
rect 4217 11396 4223 11398
rect 3915 11376 4223 11396
rect 9846 11452 10154 11472
rect 9846 11450 9852 11452
rect 9908 11450 9932 11452
rect 9988 11450 10012 11452
rect 10068 11450 10092 11452
rect 10148 11450 10154 11452
rect 9908 11398 9910 11450
rect 10090 11398 10092 11450
rect 9846 11396 9852 11398
rect 9908 11396 9932 11398
rect 9988 11396 10012 11398
rect 10068 11396 10092 11398
rect 10148 11396 10154 11398
rect 9846 11376 10154 11396
rect 6880 10908 7188 10928
rect 6880 10906 6886 10908
rect 6942 10906 6966 10908
rect 7022 10906 7046 10908
rect 7102 10906 7126 10908
rect 7182 10906 7188 10908
rect 6942 10854 6944 10906
rect 7124 10854 7126 10906
rect 6880 10852 6886 10854
rect 6942 10852 6966 10854
rect 7022 10852 7046 10854
rect 7102 10852 7126 10854
rect 7182 10852 7188 10854
rect 6880 10832 7188 10852
rect 3915 10364 4223 10384
rect 3915 10362 3921 10364
rect 3977 10362 4001 10364
rect 4057 10362 4081 10364
rect 4137 10362 4161 10364
rect 4217 10362 4223 10364
rect 3977 10310 3979 10362
rect 4159 10310 4161 10362
rect 3915 10308 3921 10310
rect 3977 10308 4001 10310
rect 4057 10308 4081 10310
rect 4137 10308 4161 10310
rect 4217 10308 4223 10310
rect 3915 10288 4223 10308
rect 9846 10364 10154 10384
rect 9846 10362 9852 10364
rect 9908 10362 9932 10364
rect 9988 10362 10012 10364
rect 10068 10362 10092 10364
rect 10148 10362 10154 10364
rect 9908 10310 9910 10362
rect 10090 10310 10092 10362
rect 9846 10308 9852 10310
rect 9908 10308 9932 10310
rect 9988 10308 10012 10310
rect 10068 10308 10092 10310
rect 10148 10308 10154 10310
rect 9846 10288 10154 10308
rect 6880 9820 7188 9840
rect 6880 9818 6886 9820
rect 6942 9818 6966 9820
rect 7022 9818 7046 9820
rect 7102 9818 7126 9820
rect 7182 9818 7188 9820
rect 6942 9766 6944 9818
rect 7124 9766 7126 9818
rect 6880 9764 6886 9766
rect 6942 9764 6966 9766
rect 7022 9764 7046 9766
rect 7102 9764 7126 9766
rect 7182 9764 7188 9766
rect 6880 9744 7188 9764
rect 3915 9276 4223 9296
rect 3915 9274 3921 9276
rect 3977 9274 4001 9276
rect 4057 9274 4081 9276
rect 4137 9274 4161 9276
rect 4217 9274 4223 9276
rect 3977 9222 3979 9274
rect 4159 9222 4161 9274
rect 3915 9220 3921 9222
rect 3977 9220 4001 9222
rect 4057 9220 4081 9222
rect 4137 9220 4161 9222
rect 4217 9220 4223 9222
rect 3915 9200 4223 9220
rect 9846 9276 10154 9296
rect 9846 9274 9852 9276
rect 9908 9274 9932 9276
rect 9988 9274 10012 9276
rect 10068 9274 10092 9276
rect 10148 9274 10154 9276
rect 9908 9222 9910 9274
rect 10090 9222 10092 9274
rect 9846 9220 9852 9222
rect 9908 9220 9932 9222
rect 9988 9220 10012 9222
rect 10068 9220 10092 9222
rect 10148 9220 10154 9222
rect 9846 9200 10154 9220
rect 6880 8732 7188 8752
rect 6880 8730 6886 8732
rect 6942 8730 6966 8732
rect 7022 8730 7046 8732
rect 7102 8730 7126 8732
rect 7182 8730 7188 8732
rect 6942 8678 6944 8730
rect 7124 8678 7126 8730
rect 6880 8676 6886 8678
rect 6942 8676 6966 8678
rect 7022 8676 7046 8678
rect 7102 8676 7126 8678
rect 7182 8676 7188 8678
rect 6880 8656 7188 8676
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1596 8265 1624 8434
rect 11348 8362 11376 17478
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1596 8090 1624 8191
rect 3915 8188 4223 8208
rect 3915 8186 3921 8188
rect 3977 8186 4001 8188
rect 4057 8186 4081 8188
rect 4137 8186 4161 8188
rect 4217 8186 4223 8188
rect 3977 8134 3979 8186
rect 4159 8134 4161 8186
rect 3915 8132 3921 8134
rect 3977 8132 4001 8134
rect 4057 8132 4081 8134
rect 4137 8132 4161 8134
rect 4217 8132 4223 8134
rect 3915 8112 4223 8132
rect 9846 8188 10154 8208
rect 9846 8186 9852 8188
rect 9908 8186 9932 8188
rect 9988 8186 10012 8188
rect 10068 8186 10092 8188
rect 10148 8186 10154 8188
rect 9908 8134 9910 8186
rect 10090 8134 10092 8186
rect 9846 8132 9852 8134
rect 9908 8132 9932 8134
rect 9988 8132 10012 8134
rect 10068 8132 10092 8134
rect 10148 8132 10154 8134
rect 9846 8112 10154 8132
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 6880 7644 7188 7664
rect 6880 7642 6886 7644
rect 6942 7642 6966 7644
rect 7022 7642 7046 7644
rect 7102 7642 7126 7644
rect 7182 7642 7188 7644
rect 6942 7590 6944 7642
rect 7124 7590 7126 7642
rect 6880 7588 6886 7590
rect 6942 7588 6966 7590
rect 7022 7588 7046 7590
rect 7102 7588 7126 7590
rect 7182 7588 7188 7590
rect 6880 7568 7188 7588
rect 3915 7100 4223 7120
rect 3915 7098 3921 7100
rect 3977 7098 4001 7100
rect 4057 7098 4081 7100
rect 4137 7098 4161 7100
rect 4217 7098 4223 7100
rect 3977 7046 3979 7098
rect 4159 7046 4161 7098
rect 3915 7044 3921 7046
rect 3977 7044 4001 7046
rect 4057 7044 4081 7046
rect 4137 7044 4161 7046
rect 4217 7044 4223 7046
rect 3915 7024 4223 7044
rect 9846 7100 10154 7120
rect 9846 7098 9852 7100
rect 9908 7098 9932 7100
rect 9988 7098 10012 7100
rect 10068 7098 10092 7100
rect 10148 7098 10154 7100
rect 9908 7046 9910 7098
rect 10090 7046 10092 7098
rect 9846 7044 9852 7046
rect 9908 7044 9932 7046
rect 9988 7044 10012 7046
rect 10068 7044 10092 7046
rect 10148 7044 10154 7046
rect 9846 7024 10154 7044
rect 6880 6556 7188 6576
rect 6880 6554 6886 6556
rect 6942 6554 6966 6556
rect 7022 6554 7046 6556
rect 7102 6554 7126 6556
rect 7182 6554 7188 6556
rect 6942 6502 6944 6554
rect 7124 6502 7126 6554
rect 6880 6500 6886 6502
rect 6942 6500 6966 6502
rect 7022 6500 7046 6502
rect 7102 6500 7126 6502
rect 7182 6500 7188 6502
rect 6880 6480 7188 6500
rect 3915 6012 4223 6032
rect 3915 6010 3921 6012
rect 3977 6010 4001 6012
rect 4057 6010 4081 6012
rect 4137 6010 4161 6012
rect 4217 6010 4223 6012
rect 3977 5958 3979 6010
rect 4159 5958 4161 6010
rect 3915 5956 3921 5958
rect 3977 5956 4001 5958
rect 4057 5956 4081 5958
rect 4137 5956 4161 5958
rect 4217 5956 4223 5958
rect 3915 5936 4223 5956
rect 9846 6012 10154 6032
rect 9846 6010 9852 6012
rect 9908 6010 9932 6012
rect 9988 6010 10012 6012
rect 10068 6010 10092 6012
rect 10148 6010 10154 6012
rect 9908 5958 9910 6010
rect 10090 5958 10092 6010
rect 9846 5956 9852 5958
rect 9908 5956 9932 5958
rect 9988 5956 10012 5958
rect 10068 5956 10092 5958
rect 10148 5956 10154 5958
rect 9846 5936 10154 5956
rect 6880 5468 7188 5488
rect 6880 5466 6886 5468
rect 6942 5466 6966 5468
rect 7022 5466 7046 5468
rect 7102 5466 7126 5468
rect 7182 5466 7188 5468
rect 6942 5414 6944 5466
rect 7124 5414 7126 5466
rect 6880 5412 6886 5414
rect 6942 5412 6966 5414
rect 7022 5412 7046 5414
rect 7102 5412 7126 5414
rect 7182 5412 7188 5414
rect 6880 5392 7188 5412
rect 3915 4924 4223 4944
rect 3915 4922 3921 4924
rect 3977 4922 4001 4924
rect 4057 4922 4081 4924
rect 4137 4922 4161 4924
rect 4217 4922 4223 4924
rect 3977 4870 3979 4922
rect 4159 4870 4161 4922
rect 3915 4868 3921 4870
rect 3977 4868 4001 4870
rect 4057 4868 4081 4870
rect 4137 4868 4161 4870
rect 4217 4868 4223 4870
rect 3915 4848 4223 4868
rect 9846 4924 10154 4944
rect 9846 4922 9852 4924
rect 9908 4922 9932 4924
rect 9988 4922 10012 4924
rect 10068 4922 10092 4924
rect 10148 4922 10154 4924
rect 9908 4870 9910 4922
rect 10090 4870 10092 4922
rect 9846 4868 9852 4870
rect 9908 4868 9932 4870
rect 9988 4868 10012 4870
rect 10068 4868 10092 4870
rect 10148 4868 10154 4870
rect 9846 4848 10154 4868
rect 6880 4380 7188 4400
rect 6880 4378 6886 4380
rect 6942 4378 6966 4380
rect 7022 4378 7046 4380
rect 7102 4378 7126 4380
rect 7182 4378 7188 4380
rect 6942 4326 6944 4378
rect 7124 4326 7126 4378
rect 6880 4324 6886 4326
rect 6942 4324 6966 4326
rect 7022 4324 7046 4326
rect 7102 4324 7126 4326
rect 7182 4324 7188 4326
rect 6880 4304 7188 4324
rect 3915 3836 4223 3856
rect 3915 3834 3921 3836
rect 3977 3834 4001 3836
rect 4057 3834 4081 3836
rect 4137 3834 4161 3836
rect 4217 3834 4223 3836
rect 3977 3782 3979 3834
rect 4159 3782 4161 3834
rect 3915 3780 3921 3782
rect 3977 3780 4001 3782
rect 4057 3780 4081 3782
rect 4137 3780 4161 3782
rect 4217 3780 4223 3782
rect 3915 3760 4223 3780
rect 9846 3836 10154 3856
rect 9846 3834 9852 3836
rect 9908 3834 9932 3836
rect 9988 3834 10012 3836
rect 10068 3834 10092 3836
rect 10148 3834 10154 3836
rect 9908 3782 9910 3834
rect 10090 3782 10092 3834
rect 9846 3780 9852 3782
rect 9908 3780 9932 3782
rect 9988 3780 10012 3782
rect 10068 3780 10092 3782
rect 10148 3780 10154 3782
rect 9846 3760 10154 3780
rect 6880 3292 7188 3312
rect 6880 3290 6886 3292
rect 6942 3290 6966 3292
rect 7022 3290 7046 3292
rect 7102 3290 7126 3292
rect 7182 3290 7188 3292
rect 6942 3238 6944 3290
rect 7124 3238 7126 3290
rect 6880 3236 6886 3238
rect 6942 3236 6966 3238
rect 7022 3236 7046 3238
rect 7102 3236 7126 3238
rect 7182 3236 7188 3238
rect 6880 3216 7188 3236
rect 2228 2984 2280 2990
rect 2226 2952 2228 2961
rect 2280 2952 2282 2961
rect 2226 2887 2282 2896
rect 1492 2848 1544 2854
rect 1490 2816 1492 2825
rect 1544 2816 1546 2825
rect 1490 2751 1546 2760
rect 3915 2748 4223 2768
rect 3915 2746 3921 2748
rect 3977 2746 4001 2748
rect 4057 2746 4081 2748
rect 4137 2746 4161 2748
rect 4217 2746 4223 2748
rect 3977 2694 3979 2746
rect 4159 2694 4161 2746
rect 3915 2692 3921 2694
rect 3977 2692 4001 2694
rect 4057 2692 4081 2694
rect 4137 2692 4161 2694
rect 4217 2692 4223 2694
rect 3915 2672 4223 2692
rect 9846 2748 10154 2768
rect 9846 2746 9852 2748
rect 9908 2746 9932 2748
rect 9988 2746 10012 2748
rect 10068 2746 10092 2748
rect 10148 2746 10154 2748
rect 9908 2694 9910 2746
rect 10090 2694 10092 2746
rect 9846 2692 9852 2694
rect 9908 2692 9932 2694
rect 9988 2692 10012 2694
rect 10068 2692 10092 2694
rect 10148 2692 10154 2694
rect 9846 2672 10154 2692
rect 12728 2650 12756 31350
rect 12811 30492 13119 30512
rect 12811 30490 12817 30492
rect 12873 30490 12897 30492
rect 12953 30490 12977 30492
rect 13033 30490 13057 30492
rect 13113 30490 13119 30492
rect 12873 30438 12875 30490
rect 13055 30438 13057 30490
rect 12811 30436 12817 30438
rect 12873 30436 12897 30438
rect 12953 30436 12977 30438
rect 13033 30436 13057 30438
rect 13113 30436 13119 30438
rect 12811 30416 13119 30436
rect 12811 29404 13119 29424
rect 12811 29402 12817 29404
rect 12873 29402 12897 29404
rect 12953 29402 12977 29404
rect 13033 29402 13057 29404
rect 13113 29402 13119 29404
rect 12873 29350 12875 29402
rect 13055 29350 13057 29402
rect 12811 29348 12817 29350
rect 12873 29348 12897 29350
rect 12953 29348 12977 29350
rect 13033 29348 13057 29350
rect 13113 29348 13119 29350
rect 12811 29328 13119 29348
rect 12811 28316 13119 28336
rect 12811 28314 12817 28316
rect 12873 28314 12897 28316
rect 12953 28314 12977 28316
rect 13033 28314 13057 28316
rect 13113 28314 13119 28316
rect 12873 28262 12875 28314
rect 13055 28262 13057 28314
rect 12811 28260 12817 28262
rect 12873 28260 12897 28262
rect 12953 28260 12977 28262
rect 13033 28260 13057 28262
rect 13113 28260 13119 28262
rect 12811 28240 13119 28260
rect 12811 27228 13119 27248
rect 12811 27226 12817 27228
rect 12873 27226 12897 27228
rect 12953 27226 12977 27228
rect 13033 27226 13057 27228
rect 13113 27226 13119 27228
rect 12873 27174 12875 27226
rect 13055 27174 13057 27226
rect 12811 27172 12817 27174
rect 12873 27172 12897 27174
rect 12953 27172 12977 27174
rect 13033 27172 13057 27174
rect 13113 27172 13119 27174
rect 12811 27152 13119 27172
rect 12811 26140 13119 26160
rect 12811 26138 12817 26140
rect 12873 26138 12897 26140
rect 12953 26138 12977 26140
rect 13033 26138 13057 26140
rect 13113 26138 13119 26140
rect 12873 26086 12875 26138
rect 13055 26086 13057 26138
rect 12811 26084 12817 26086
rect 12873 26084 12897 26086
rect 12953 26084 12977 26086
rect 13033 26084 13057 26086
rect 13113 26084 13119 26086
rect 12811 26064 13119 26084
rect 13174 25528 13230 25537
rect 13174 25463 13176 25472
rect 13228 25463 13230 25472
rect 13176 25434 13228 25440
rect 12811 25052 13119 25072
rect 12811 25050 12817 25052
rect 12873 25050 12897 25052
rect 12953 25050 12977 25052
rect 13033 25050 13057 25052
rect 13113 25050 13119 25052
rect 12873 24998 12875 25050
rect 13055 24998 13057 25050
rect 12811 24996 12817 24998
rect 12873 24996 12897 24998
rect 12953 24996 12977 24998
rect 13033 24996 13057 24998
rect 13113 24996 13119 24998
rect 12811 24976 13119 24996
rect 13188 24886 13216 25434
rect 13176 24880 13228 24886
rect 13176 24822 13228 24828
rect 13188 24342 13216 24822
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 13188 24206 13216 24278
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 12811 23964 13119 23984
rect 12811 23962 12817 23964
rect 12873 23962 12897 23964
rect 12953 23962 12977 23964
rect 13033 23962 13057 23964
rect 13113 23962 13119 23964
rect 12873 23910 12875 23962
rect 13055 23910 13057 23962
rect 12811 23908 12817 23910
rect 12873 23908 12897 23910
rect 12953 23908 12977 23910
rect 13033 23908 13057 23910
rect 13113 23908 13119 23910
rect 12811 23888 13119 23908
rect 12811 22876 13119 22896
rect 12811 22874 12817 22876
rect 12873 22874 12897 22876
rect 12953 22874 12977 22876
rect 13033 22874 13057 22876
rect 13113 22874 13119 22876
rect 12873 22822 12875 22874
rect 13055 22822 13057 22874
rect 12811 22820 12817 22822
rect 12873 22820 12897 22822
rect 12953 22820 12977 22822
rect 13033 22820 13057 22822
rect 13113 22820 13119 22822
rect 12811 22800 13119 22820
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 12811 21788 13119 21808
rect 12811 21786 12817 21788
rect 12873 21786 12897 21788
rect 12953 21786 12977 21788
rect 13033 21786 13057 21788
rect 13113 21786 13119 21788
rect 12873 21734 12875 21786
rect 13055 21734 13057 21786
rect 12811 21732 12817 21734
rect 12873 21732 12897 21734
rect 12953 21732 12977 21734
rect 13033 21732 13057 21734
rect 13113 21732 13119 21734
rect 12811 21712 13119 21732
rect 12811 20700 13119 20720
rect 12811 20698 12817 20700
rect 12873 20698 12897 20700
rect 12953 20698 12977 20700
rect 13033 20698 13057 20700
rect 13113 20698 13119 20700
rect 12873 20646 12875 20698
rect 13055 20646 13057 20698
rect 12811 20644 12817 20646
rect 12873 20644 12897 20646
rect 12953 20644 12977 20646
rect 13033 20644 13057 20646
rect 13113 20644 13119 20646
rect 12811 20624 13119 20644
rect 13280 20466 13308 21830
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 12811 19612 13119 19632
rect 12811 19610 12817 19612
rect 12873 19610 12897 19612
rect 12953 19610 12977 19612
rect 13033 19610 13057 19612
rect 13113 19610 13119 19612
rect 12873 19558 12875 19610
rect 13055 19558 13057 19610
rect 12811 19556 12817 19558
rect 12873 19556 12897 19558
rect 12953 19556 12977 19558
rect 13033 19556 13057 19558
rect 13113 19556 13119 19558
rect 12811 19536 13119 19556
rect 12811 18524 13119 18544
rect 12811 18522 12817 18524
rect 12873 18522 12897 18524
rect 12953 18522 12977 18524
rect 13033 18522 13057 18524
rect 13113 18522 13119 18524
rect 12873 18470 12875 18522
rect 13055 18470 13057 18522
rect 12811 18468 12817 18470
rect 12873 18468 12897 18470
rect 12953 18468 12977 18470
rect 13033 18468 13057 18470
rect 13113 18468 13119 18470
rect 12811 18448 13119 18468
rect 13280 18358 13308 20402
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 12811 17436 13119 17456
rect 12811 17434 12817 17436
rect 12873 17434 12897 17436
rect 12953 17434 12977 17436
rect 13033 17434 13057 17436
rect 13113 17434 13119 17436
rect 12873 17382 12875 17434
rect 13055 17382 13057 17434
rect 12811 17380 12817 17382
rect 12873 17380 12897 17382
rect 12953 17380 12977 17382
rect 13033 17380 13057 17382
rect 13113 17380 13119 17382
rect 12811 17360 13119 17380
rect 12811 16348 13119 16368
rect 12811 16346 12817 16348
rect 12873 16346 12897 16348
rect 12953 16346 12977 16348
rect 13033 16346 13057 16348
rect 13113 16346 13119 16348
rect 12873 16294 12875 16346
rect 13055 16294 13057 16346
rect 12811 16292 12817 16294
rect 12873 16292 12897 16294
rect 12953 16292 12977 16294
rect 13033 16292 13057 16294
rect 13113 16292 13119 16294
rect 12811 16272 13119 16292
rect 12811 15260 13119 15280
rect 12811 15258 12817 15260
rect 12873 15258 12897 15260
rect 12953 15258 12977 15260
rect 13033 15258 13057 15260
rect 13113 15258 13119 15260
rect 12873 15206 12875 15258
rect 13055 15206 13057 15258
rect 12811 15204 12817 15206
rect 12873 15204 12897 15206
rect 12953 15204 12977 15206
rect 13033 15204 13057 15206
rect 13113 15204 13119 15206
rect 12811 15184 13119 15204
rect 12811 14172 13119 14192
rect 12811 14170 12817 14172
rect 12873 14170 12897 14172
rect 12953 14170 12977 14172
rect 13033 14170 13057 14172
rect 13113 14170 13119 14172
rect 12873 14118 12875 14170
rect 13055 14118 13057 14170
rect 12811 14116 12817 14118
rect 12873 14116 12897 14118
rect 12953 14116 12977 14118
rect 13033 14116 13057 14118
rect 13113 14116 13119 14118
rect 12811 14096 13119 14116
rect 12811 13084 13119 13104
rect 12811 13082 12817 13084
rect 12873 13082 12897 13084
rect 12953 13082 12977 13084
rect 13033 13082 13057 13084
rect 13113 13082 13119 13084
rect 12873 13030 12875 13082
rect 13055 13030 13057 13082
rect 12811 13028 12817 13030
rect 12873 13028 12897 13030
rect 12953 13028 12977 13030
rect 13033 13028 13057 13030
rect 13113 13028 13119 13030
rect 12811 13008 13119 13028
rect 12811 11996 13119 12016
rect 12811 11994 12817 11996
rect 12873 11994 12897 11996
rect 12953 11994 12977 11996
rect 13033 11994 13057 11996
rect 13113 11994 13119 11996
rect 12873 11942 12875 11994
rect 13055 11942 13057 11994
rect 12811 11940 12817 11942
rect 12873 11940 12897 11942
rect 12953 11940 12977 11942
rect 13033 11940 13057 11942
rect 13113 11940 13119 11942
rect 12811 11920 13119 11940
rect 12811 10908 13119 10928
rect 12811 10906 12817 10908
rect 12873 10906 12897 10908
rect 12953 10906 12977 10908
rect 13033 10906 13057 10908
rect 13113 10906 13119 10908
rect 12873 10854 12875 10906
rect 13055 10854 13057 10906
rect 12811 10852 12817 10854
rect 12873 10852 12897 10854
rect 12953 10852 12977 10854
rect 13033 10852 13057 10854
rect 13113 10852 13119 10854
rect 12811 10832 13119 10852
rect 12811 9820 13119 9840
rect 12811 9818 12817 9820
rect 12873 9818 12897 9820
rect 12953 9818 12977 9820
rect 13033 9818 13057 9820
rect 13113 9818 13119 9820
rect 12873 9766 12875 9818
rect 13055 9766 13057 9818
rect 12811 9764 12817 9766
rect 12873 9764 12897 9766
rect 12953 9764 12977 9766
rect 13033 9764 13057 9766
rect 13113 9764 13119 9766
rect 12811 9744 13119 9764
rect 12811 8732 13119 8752
rect 12811 8730 12817 8732
rect 12873 8730 12897 8732
rect 12953 8730 12977 8732
rect 13033 8730 13057 8732
rect 13113 8730 13119 8732
rect 12873 8678 12875 8730
rect 13055 8678 13057 8730
rect 12811 8676 12817 8678
rect 12873 8676 12897 8678
rect 12953 8676 12977 8678
rect 13033 8676 13057 8678
rect 13113 8676 13119 8678
rect 12811 8656 13119 8676
rect 12811 7644 13119 7664
rect 12811 7642 12817 7644
rect 12873 7642 12897 7644
rect 12953 7642 12977 7644
rect 13033 7642 13057 7644
rect 13113 7642 13119 7644
rect 12873 7590 12875 7642
rect 13055 7590 13057 7642
rect 12811 7588 12817 7590
rect 12873 7588 12897 7590
rect 12953 7588 12977 7590
rect 13033 7588 13057 7590
rect 13113 7588 13119 7590
rect 12811 7568 13119 7588
rect 12811 6556 13119 6576
rect 12811 6554 12817 6556
rect 12873 6554 12897 6556
rect 12953 6554 12977 6556
rect 13033 6554 13057 6556
rect 13113 6554 13119 6556
rect 12873 6502 12875 6554
rect 13055 6502 13057 6554
rect 12811 6500 12817 6502
rect 12873 6500 12897 6502
rect 12953 6500 12977 6502
rect 13033 6500 13057 6502
rect 13113 6500 13119 6502
rect 12811 6480 13119 6500
rect 12811 5468 13119 5488
rect 12811 5466 12817 5468
rect 12873 5466 12897 5468
rect 12953 5466 12977 5468
rect 13033 5466 13057 5468
rect 13113 5466 13119 5468
rect 12873 5414 12875 5466
rect 13055 5414 13057 5466
rect 12811 5412 12817 5414
rect 12873 5412 12897 5414
rect 12953 5412 12977 5414
rect 13033 5412 13057 5414
rect 13113 5412 13119 5414
rect 12811 5392 13119 5412
rect 12811 4380 13119 4400
rect 12811 4378 12817 4380
rect 12873 4378 12897 4380
rect 12953 4378 12977 4380
rect 13033 4378 13057 4380
rect 13113 4378 13119 4380
rect 12873 4326 12875 4378
rect 13055 4326 13057 4378
rect 12811 4324 12817 4326
rect 12873 4324 12897 4326
rect 12953 4324 12977 4326
rect 13033 4324 13057 4326
rect 13113 4324 13119 4326
rect 12811 4304 13119 4324
rect 12811 3292 13119 3312
rect 12811 3290 12817 3292
rect 12873 3290 12897 3292
rect 12953 3290 12977 3292
rect 13033 3290 13057 3292
rect 13113 3290 13119 3292
rect 12873 3238 12875 3290
rect 13055 3238 13057 3290
rect 12811 3236 12817 3238
rect 12873 3236 12897 3238
rect 12953 3236 12977 3238
rect 13033 3236 13057 3238
rect 13113 3236 13119 3238
rect 12811 3216 13119 3236
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 2504 2372 2556 2378
rect 2504 2314 2556 2320
rect 2516 800 2544 2314
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 6880 2204 7188 2224
rect 6880 2202 6886 2204
rect 6942 2202 6966 2204
rect 7022 2202 7046 2204
rect 7102 2202 7126 2204
rect 7182 2202 7188 2204
rect 6942 2150 6944 2202
rect 7124 2150 7126 2202
rect 6880 2148 6886 2150
rect 6942 2148 6966 2150
rect 7022 2148 7046 2150
rect 7102 2148 7126 2150
rect 7182 2148 7188 2150
rect 6880 2128 7188 2148
rect 7484 800 7512 2246
rect 12452 800 12480 2382
rect 13372 2378 13400 31758
rect 13648 29510 13676 32506
rect 13636 29504 13688 29510
rect 13636 29446 13688 29452
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13452 25832 13504 25838
rect 13452 25774 13504 25780
rect 13464 24818 13492 25774
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13464 24410 13492 24754
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13556 24274 13584 24550
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13648 24138 13676 25842
rect 13636 24132 13688 24138
rect 13636 24074 13688 24080
rect 13648 22098 13676 24074
rect 14016 22098 14044 47126
rect 14200 46714 14228 49286
rect 14554 49286 14780 49314
rect 14554 49200 14610 49286
rect 14188 46708 14240 46714
rect 14188 46650 14240 46656
rect 14752 46170 14780 49286
rect 14844 49286 15070 49314
rect 14844 47054 14872 49286
rect 15014 49200 15070 49286
rect 15474 49200 15530 50000
rect 15934 49314 15990 50000
rect 16394 49314 16450 50000
rect 16854 49314 16910 50000
rect 17314 49314 17370 50000
rect 15934 49286 16160 49314
rect 15934 49200 15990 49286
rect 14832 47048 14884 47054
rect 14832 46990 14884 46996
rect 15292 47048 15344 47054
rect 15292 46990 15344 46996
rect 15108 46572 15160 46578
rect 15108 46514 15160 46520
rect 14740 46164 14792 46170
rect 14740 46106 14792 46112
rect 14280 36032 14332 36038
rect 14280 35974 14332 35980
rect 14292 33590 14320 35974
rect 15120 35562 15148 46514
rect 15200 36236 15252 36242
rect 15200 36178 15252 36184
rect 15108 35556 15160 35562
rect 15108 35498 15160 35504
rect 14464 35488 14516 35494
rect 14464 35430 14516 35436
rect 14372 35216 14424 35222
rect 14372 35158 14424 35164
rect 14384 34610 14412 35158
rect 14476 34678 14504 35430
rect 14832 35148 14884 35154
rect 14832 35090 14884 35096
rect 14464 34672 14516 34678
rect 14464 34614 14516 34620
rect 14372 34604 14424 34610
rect 14372 34546 14424 34552
rect 14476 33998 14504 34614
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14648 33924 14700 33930
rect 14648 33866 14700 33872
rect 14280 33584 14332 33590
rect 14280 33526 14332 33532
rect 14292 32910 14320 33526
rect 14660 33522 14688 33866
rect 14752 33658 14780 34546
rect 14844 34474 14872 35090
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 14924 35012 14976 35018
rect 14924 34954 14976 34960
rect 14936 34610 14964 34954
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 14832 34468 14884 34474
rect 14832 34410 14884 34416
rect 14924 33856 14976 33862
rect 14924 33798 14976 33804
rect 14936 33658 14964 33798
rect 14740 33652 14792 33658
rect 14740 33594 14792 33600
rect 14924 33652 14976 33658
rect 14924 33594 14976 33600
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14648 33516 14700 33522
rect 14648 33458 14700 33464
rect 14568 32978 14596 33458
rect 15028 33454 15056 34546
rect 15120 33862 15148 35022
rect 15212 34746 15240 36178
rect 15200 34740 15252 34746
rect 15200 34682 15252 34688
rect 15108 33856 15160 33862
rect 15108 33798 15160 33804
rect 15016 33448 15068 33454
rect 15016 33390 15068 33396
rect 14740 33312 14792 33318
rect 14740 33254 14792 33260
rect 14752 33046 14780 33254
rect 15120 33114 15148 33798
rect 15200 33584 15252 33590
rect 15200 33526 15252 33532
rect 15212 33318 15240 33526
rect 15200 33312 15252 33318
rect 15200 33254 15252 33260
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 14740 33040 14792 33046
rect 14740 32982 14792 32988
rect 14556 32972 14608 32978
rect 14556 32914 14608 32920
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 14752 32434 14780 32982
rect 15200 32904 15252 32910
rect 15200 32846 15252 32852
rect 14832 32836 14884 32842
rect 14832 32778 14884 32784
rect 14844 32434 14872 32778
rect 15212 32570 15240 32846
rect 15200 32564 15252 32570
rect 15200 32506 15252 32512
rect 15304 32502 15332 46990
rect 15488 46646 15516 49200
rect 15776 47356 16084 47376
rect 15776 47354 15782 47356
rect 15838 47354 15862 47356
rect 15918 47354 15942 47356
rect 15998 47354 16022 47356
rect 16078 47354 16084 47356
rect 15838 47302 15840 47354
rect 16020 47302 16022 47354
rect 15776 47300 15782 47302
rect 15838 47300 15862 47302
rect 15918 47300 15942 47302
rect 15998 47300 16022 47302
rect 16078 47300 16084 47302
rect 15776 47280 16084 47300
rect 16132 47122 16160 49286
rect 16394 49286 16528 49314
rect 16394 49200 16450 49286
rect 16500 47122 16528 49286
rect 16854 49286 16988 49314
rect 16854 49200 16910 49286
rect 16120 47116 16172 47122
rect 16120 47058 16172 47064
rect 16488 47116 16540 47122
rect 16488 47058 16540 47064
rect 16132 46714 16160 47058
rect 16856 47048 16908 47054
rect 16486 47016 16542 47025
rect 16856 46990 16908 46996
rect 16486 46951 16542 46960
rect 16120 46708 16172 46714
rect 16120 46650 16172 46656
rect 15476 46640 15528 46646
rect 15476 46582 15528 46588
rect 15488 46170 15516 46582
rect 15660 46572 15712 46578
rect 15660 46514 15712 46520
rect 15568 46436 15620 46442
rect 15568 46378 15620 46384
rect 15476 46164 15528 46170
rect 15476 46106 15528 46112
rect 15580 45937 15608 46378
rect 15566 45928 15622 45937
rect 15566 45863 15622 45872
rect 15672 45554 15700 46514
rect 15776 46268 16084 46288
rect 15776 46266 15782 46268
rect 15838 46266 15862 46268
rect 15918 46266 15942 46268
rect 15998 46266 16022 46268
rect 16078 46266 16084 46268
rect 15838 46214 15840 46266
rect 16020 46214 16022 46266
rect 15776 46212 15782 46214
rect 15838 46212 15862 46214
rect 15918 46212 15942 46214
rect 15998 46212 16022 46214
rect 16078 46212 16084 46214
rect 15776 46192 16084 46212
rect 15580 45526 15700 45554
rect 15476 44804 15528 44810
rect 15476 44746 15528 44752
rect 15488 34746 15516 44746
rect 15580 35766 15608 45526
rect 15776 45180 16084 45200
rect 15776 45178 15782 45180
rect 15838 45178 15862 45180
rect 15918 45178 15942 45180
rect 15998 45178 16022 45180
rect 16078 45178 16084 45180
rect 15838 45126 15840 45178
rect 16020 45126 16022 45178
rect 15776 45124 15782 45126
rect 15838 45124 15862 45126
rect 15918 45124 15942 45126
rect 15998 45124 16022 45126
rect 16078 45124 16084 45126
rect 15776 45104 16084 45124
rect 16500 44538 16528 46951
rect 16488 44532 16540 44538
rect 16488 44474 16540 44480
rect 15776 44092 16084 44112
rect 15776 44090 15782 44092
rect 15838 44090 15862 44092
rect 15918 44090 15942 44092
rect 15998 44090 16022 44092
rect 16078 44090 16084 44092
rect 15838 44038 15840 44090
rect 16020 44038 16022 44090
rect 15776 44036 15782 44038
rect 15838 44036 15862 44038
rect 15918 44036 15942 44038
rect 15998 44036 16022 44038
rect 16078 44036 16084 44038
rect 15776 44016 16084 44036
rect 15776 43004 16084 43024
rect 15776 43002 15782 43004
rect 15838 43002 15862 43004
rect 15918 43002 15942 43004
rect 15998 43002 16022 43004
rect 16078 43002 16084 43004
rect 15838 42950 15840 43002
rect 16020 42950 16022 43002
rect 15776 42948 15782 42950
rect 15838 42948 15862 42950
rect 15918 42948 15942 42950
rect 15998 42948 16022 42950
rect 16078 42948 16084 42950
rect 15776 42928 16084 42948
rect 15776 41916 16084 41936
rect 15776 41914 15782 41916
rect 15838 41914 15862 41916
rect 15918 41914 15942 41916
rect 15998 41914 16022 41916
rect 16078 41914 16084 41916
rect 15838 41862 15840 41914
rect 16020 41862 16022 41914
rect 15776 41860 15782 41862
rect 15838 41860 15862 41862
rect 15918 41860 15942 41862
rect 15998 41860 16022 41862
rect 16078 41860 16084 41862
rect 15776 41840 16084 41860
rect 15776 40828 16084 40848
rect 15776 40826 15782 40828
rect 15838 40826 15862 40828
rect 15918 40826 15942 40828
rect 15998 40826 16022 40828
rect 16078 40826 16084 40828
rect 15838 40774 15840 40826
rect 16020 40774 16022 40826
rect 15776 40772 15782 40774
rect 15838 40772 15862 40774
rect 15918 40772 15942 40774
rect 15998 40772 16022 40774
rect 16078 40772 16084 40774
rect 15776 40752 16084 40772
rect 15776 39740 16084 39760
rect 15776 39738 15782 39740
rect 15838 39738 15862 39740
rect 15918 39738 15942 39740
rect 15998 39738 16022 39740
rect 16078 39738 16084 39740
rect 15838 39686 15840 39738
rect 16020 39686 16022 39738
rect 15776 39684 15782 39686
rect 15838 39684 15862 39686
rect 15918 39684 15942 39686
rect 15998 39684 16022 39686
rect 16078 39684 16084 39686
rect 15776 39664 16084 39684
rect 15776 38652 16084 38672
rect 15776 38650 15782 38652
rect 15838 38650 15862 38652
rect 15918 38650 15942 38652
rect 15998 38650 16022 38652
rect 16078 38650 16084 38652
rect 15838 38598 15840 38650
rect 16020 38598 16022 38650
rect 15776 38596 15782 38598
rect 15838 38596 15862 38598
rect 15918 38596 15942 38598
rect 15998 38596 16022 38598
rect 16078 38596 16084 38598
rect 15776 38576 16084 38596
rect 15776 37564 16084 37584
rect 15776 37562 15782 37564
rect 15838 37562 15862 37564
rect 15918 37562 15942 37564
rect 15998 37562 16022 37564
rect 16078 37562 16084 37564
rect 15838 37510 15840 37562
rect 16020 37510 16022 37562
rect 15776 37508 15782 37510
rect 15838 37508 15862 37510
rect 15918 37508 15942 37510
rect 15998 37508 16022 37510
rect 16078 37508 16084 37510
rect 15776 37488 16084 37508
rect 16396 37188 16448 37194
rect 16396 37130 16448 37136
rect 15776 36476 16084 36496
rect 15776 36474 15782 36476
rect 15838 36474 15862 36476
rect 15918 36474 15942 36476
rect 15998 36474 16022 36476
rect 16078 36474 16084 36476
rect 15838 36422 15840 36474
rect 16020 36422 16022 36474
rect 15776 36420 15782 36422
rect 15838 36420 15862 36422
rect 15918 36420 15942 36422
rect 15998 36420 16022 36422
rect 16078 36420 16084 36422
rect 15776 36400 16084 36420
rect 15660 36032 15712 36038
rect 15660 35974 15712 35980
rect 16304 36032 16356 36038
rect 16304 35974 16356 35980
rect 15568 35760 15620 35766
rect 15568 35702 15620 35708
rect 15476 34740 15528 34746
rect 15476 34682 15528 34688
rect 15384 34536 15436 34542
rect 15384 34478 15436 34484
rect 15292 32496 15344 32502
rect 15292 32438 15344 32444
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14740 32428 14792 32434
rect 14740 32370 14792 32376
rect 14832 32428 14884 32434
rect 14832 32370 14884 32376
rect 14108 31346 14136 32370
rect 15016 32224 15068 32230
rect 15016 32166 15068 32172
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15028 32026 15056 32166
rect 15016 32020 15068 32026
rect 15016 31962 15068 31968
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 14096 31340 14148 31346
rect 14096 31282 14148 31288
rect 14108 30734 14136 31282
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 14372 29708 14424 29714
rect 14372 29650 14424 29656
rect 14384 26042 14412 29650
rect 14372 26036 14424 26042
rect 14372 25978 14424 25984
rect 14188 25832 14240 25838
rect 14188 25774 14240 25780
rect 14200 24818 14228 25774
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 13452 22024 13504 22030
rect 13452 21966 13504 21972
rect 13464 20466 13492 21966
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13464 18426 13492 20402
rect 14016 19310 14044 22034
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 14752 2582 14780 31826
rect 15212 30870 15240 32166
rect 15304 31278 15332 32438
rect 15292 31272 15344 31278
rect 15292 31214 15344 31220
rect 15200 30864 15252 30870
rect 15200 30806 15252 30812
rect 15396 30326 15424 34478
rect 15488 33998 15516 34682
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15488 33810 15516 33934
rect 15580 33930 15608 35702
rect 15672 35698 15700 35974
rect 15660 35692 15712 35698
rect 15660 35634 15712 35640
rect 15672 34513 15700 35634
rect 16212 35624 16264 35630
rect 16212 35566 16264 35572
rect 15776 35388 16084 35408
rect 15776 35386 15782 35388
rect 15838 35386 15862 35388
rect 15918 35386 15942 35388
rect 15998 35386 16022 35388
rect 16078 35386 16084 35388
rect 15838 35334 15840 35386
rect 16020 35334 16022 35386
rect 15776 35332 15782 35334
rect 15838 35332 15862 35334
rect 15918 35332 15942 35334
rect 15998 35332 16022 35334
rect 16078 35332 16084 35334
rect 15776 35312 16084 35332
rect 16028 35216 16080 35222
rect 16028 35158 16080 35164
rect 16040 34950 16068 35158
rect 16028 34944 16080 34950
rect 16028 34886 16080 34892
rect 15750 34640 15806 34649
rect 15750 34575 15806 34584
rect 15658 34504 15714 34513
rect 15658 34439 15714 34448
rect 15764 34388 15792 34575
rect 15672 34360 15792 34388
rect 15672 34066 15700 34360
rect 15776 34300 16084 34320
rect 15776 34298 15782 34300
rect 15838 34298 15862 34300
rect 15918 34298 15942 34300
rect 15998 34298 16022 34300
rect 16078 34298 16084 34300
rect 15838 34246 15840 34298
rect 16020 34246 16022 34298
rect 15776 34244 15782 34246
rect 15838 34244 15862 34246
rect 15918 34244 15942 34246
rect 15998 34244 16022 34246
rect 16078 34244 16084 34246
rect 15776 34224 16084 34244
rect 15660 34060 15712 34066
rect 15660 34002 15712 34008
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 15568 33924 15620 33930
rect 15568 33866 15620 33872
rect 15488 33782 15884 33810
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 15580 33561 15608 33594
rect 15566 33552 15622 33561
rect 15856 33522 15884 33782
rect 16040 33590 16068 33934
rect 16028 33584 16080 33590
rect 16028 33526 16080 33532
rect 15566 33487 15622 33496
rect 15844 33516 15896 33522
rect 15844 33458 15896 33464
rect 16224 33454 16252 35566
rect 16212 33448 16264 33454
rect 16212 33390 16264 33396
rect 15776 33212 16084 33232
rect 15776 33210 15782 33212
rect 15838 33210 15862 33212
rect 15918 33210 15942 33212
rect 15998 33210 16022 33212
rect 16078 33210 16084 33212
rect 15838 33158 15840 33210
rect 16020 33158 16022 33210
rect 15776 33156 15782 33158
rect 15838 33156 15862 33158
rect 15918 33156 15942 33158
rect 15998 33156 16022 33158
rect 16078 33156 16084 33158
rect 15776 33136 16084 33156
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 15476 32020 15528 32026
rect 15476 31962 15528 31968
rect 15488 30734 15516 31962
rect 15580 31482 15608 32370
rect 16040 32298 16160 32314
rect 16028 32292 16160 32298
rect 16080 32286 16160 32292
rect 16028 32234 16080 32240
rect 15776 32124 16084 32144
rect 15776 32122 15782 32124
rect 15838 32122 15862 32124
rect 15918 32122 15942 32124
rect 15998 32122 16022 32124
rect 16078 32122 16084 32124
rect 15838 32070 15840 32122
rect 16020 32070 16022 32122
rect 15776 32068 15782 32070
rect 15838 32068 15862 32070
rect 15918 32068 15942 32070
rect 15998 32068 16022 32070
rect 16078 32068 16084 32070
rect 15776 32048 16084 32068
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 16132 31210 16160 32286
rect 16120 31204 16172 31210
rect 16120 31146 16172 31152
rect 15776 31036 16084 31056
rect 15776 31034 15782 31036
rect 15838 31034 15862 31036
rect 15918 31034 15942 31036
rect 15998 31034 16022 31036
rect 16078 31034 16084 31036
rect 15838 30982 15840 31034
rect 16020 30982 16022 31034
rect 15776 30980 15782 30982
rect 15838 30980 15862 30982
rect 15918 30980 15942 30982
rect 15998 30980 16022 30982
rect 16078 30980 16084 30982
rect 15776 30960 16084 30980
rect 16132 30818 16160 31146
rect 16040 30790 16160 30818
rect 16040 30734 16068 30790
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 16028 30728 16080 30734
rect 16028 30670 16080 30676
rect 15752 30592 15804 30598
rect 15752 30534 15804 30540
rect 15384 30320 15436 30326
rect 15384 30262 15436 30268
rect 15764 30258 15792 30534
rect 16040 30258 16068 30670
rect 15752 30252 15804 30258
rect 15752 30194 15804 30200
rect 16028 30252 16080 30258
rect 16028 30194 16080 30200
rect 15108 30184 15160 30190
rect 15764 30138 15792 30194
rect 15108 30126 15160 30132
rect 15120 29714 15148 30126
rect 15672 30110 15792 30138
rect 15108 29708 15160 29714
rect 15108 29650 15160 29656
rect 15672 29646 15700 30110
rect 15776 29948 16084 29968
rect 15776 29946 15782 29948
rect 15838 29946 15862 29948
rect 15918 29946 15942 29948
rect 15998 29946 16022 29948
rect 16078 29946 16084 29948
rect 15838 29894 15840 29946
rect 16020 29894 16022 29946
rect 15776 29892 15782 29894
rect 15838 29892 15862 29894
rect 15918 29892 15942 29894
rect 15998 29892 16022 29894
rect 16078 29892 16084 29894
rect 15776 29872 16084 29892
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15568 29504 15620 29510
rect 15568 29446 15620 29452
rect 15580 26234 15608 29446
rect 15776 28860 16084 28880
rect 15776 28858 15782 28860
rect 15838 28858 15862 28860
rect 15918 28858 15942 28860
rect 15998 28858 16022 28860
rect 16078 28858 16084 28860
rect 15838 28806 15840 28858
rect 16020 28806 16022 28858
rect 15776 28804 15782 28806
rect 15838 28804 15862 28806
rect 15918 28804 15942 28806
rect 15998 28804 16022 28806
rect 16078 28804 16084 28806
rect 15776 28784 16084 28804
rect 16224 28762 16252 33390
rect 16316 33318 16344 35974
rect 16408 34610 16436 37130
rect 16868 36174 16896 46990
rect 16960 46034 16988 49286
rect 17314 49286 17448 49314
rect 17314 49200 17370 49286
rect 17316 46504 17368 46510
rect 17316 46446 17368 46452
rect 16948 46028 17000 46034
rect 16948 45970 17000 45976
rect 16960 45082 16988 45970
rect 17040 45960 17092 45966
rect 17040 45902 17092 45908
rect 17224 45960 17276 45966
rect 17224 45902 17276 45908
rect 16948 45076 17000 45082
rect 16948 45018 17000 45024
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16580 36100 16632 36106
rect 16580 36042 16632 36048
rect 16592 35698 16620 36042
rect 16868 35698 16896 36110
rect 16580 35692 16632 35698
rect 16580 35634 16632 35640
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16856 35488 16908 35494
rect 16856 35430 16908 35436
rect 16580 35080 16632 35086
rect 16580 35022 16632 35028
rect 16396 34604 16448 34610
rect 16396 34546 16448 34552
rect 16408 34066 16436 34546
rect 16488 34536 16540 34542
rect 16488 34478 16540 34484
rect 16500 34202 16528 34478
rect 16592 34406 16620 35022
rect 16764 34604 16816 34610
rect 16764 34546 16816 34552
rect 16580 34400 16632 34406
rect 16580 34342 16632 34348
rect 16488 34196 16540 34202
rect 16488 34138 16540 34144
rect 16396 34060 16448 34066
rect 16396 34002 16448 34008
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16304 33312 16356 33318
rect 16592 33289 16620 33866
rect 16304 33254 16356 33260
rect 16578 33280 16634 33289
rect 16316 32910 16344 33254
rect 16578 33215 16634 33224
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16316 31754 16344 32846
rect 16592 32434 16620 33050
rect 16580 32428 16632 32434
rect 16580 32370 16632 32376
rect 16684 32298 16712 33934
rect 16776 33590 16804 34546
rect 16764 33584 16816 33590
rect 16764 33526 16816 33532
rect 16868 33386 16896 35430
rect 16960 34649 16988 37062
rect 17052 36922 17080 45902
rect 17132 45484 17184 45490
rect 17132 45426 17184 45432
rect 17040 36916 17092 36922
rect 17040 36858 17092 36864
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 16946 34640 17002 34649
rect 16946 34575 16948 34584
rect 17000 34575 17002 34584
rect 16948 34546 17000 34552
rect 16960 34515 16988 34546
rect 16948 34400 17000 34406
rect 16948 34342 17000 34348
rect 16960 33522 16988 34342
rect 17052 33998 17080 35634
rect 17144 34474 17172 45426
rect 17236 36106 17264 45902
rect 17328 45558 17356 46446
rect 17316 45552 17368 45558
rect 17316 45494 17368 45500
rect 17420 45354 17448 49286
rect 17774 49200 17830 50000
rect 18234 49314 18290 50000
rect 18694 49314 18750 50000
rect 18234 49286 18368 49314
rect 18234 49200 18290 49286
rect 17788 46170 17816 49200
rect 18236 47456 18288 47462
rect 18236 47398 18288 47404
rect 17776 46164 17828 46170
rect 17776 46106 17828 46112
rect 18052 45484 18104 45490
rect 18052 45426 18104 45432
rect 17408 45348 17460 45354
rect 17408 45290 17460 45296
rect 17592 45348 17644 45354
rect 17592 45290 17644 45296
rect 17224 36100 17276 36106
rect 17224 36042 17276 36048
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17132 34468 17184 34474
rect 17132 34410 17184 34416
rect 17512 34066 17540 35226
rect 17500 34060 17552 34066
rect 17500 34002 17552 34008
rect 17040 33992 17092 33998
rect 17040 33934 17092 33940
rect 17604 33561 17632 45290
rect 18064 45082 18092 45426
rect 18052 45076 18104 45082
rect 18052 45018 18104 45024
rect 18248 44878 18276 47398
rect 18340 45490 18368 49286
rect 18432 49286 18750 49314
rect 18432 47462 18460 49286
rect 18694 49200 18750 49286
rect 19154 49200 19210 50000
rect 19614 49200 19670 50000
rect 18420 47456 18472 47462
rect 18420 47398 18472 47404
rect 19168 46646 19196 49200
rect 19156 46640 19208 46646
rect 19156 46582 19208 46588
rect 19628 46510 19656 49200
rect 19616 46504 19668 46510
rect 19616 46446 19668 46452
rect 18328 45484 18380 45490
rect 18328 45426 18380 45432
rect 18236 44872 18288 44878
rect 18236 44814 18288 44820
rect 18248 44470 18276 44814
rect 18236 44464 18288 44470
rect 18236 44406 18288 44412
rect 18052 44396 18104 44402
rect 18052 44338 18104 44344
rect 17960 40928 18012 40934
rect 17960 40870 18012 40876
rect 17972 37262 18000 40870
rect 17960 37256 18012 37262
rect 17960 37198 18012 37204
rect 17972 36854 18000 37198
rect 17960 36848 18012 36854
rect 17960 36790 18012 36796
rect 17776 36576 17828 36582
rect 17776 36518 17828 36524
rect 17788 34950 17816 36518
rect 18064 36378 18092 44338
rect 18144 41132 18196 41138
rect 18144 41074 18196 41080
rect 18156 40769 18184 41074
rect 18142 40760 18198 40769
rect 18142 40695 18198 40704
rect 18144 37256 18196 37262
rect 18144 37198 18196 37204
rect 18156 36786 18184 37198
rect 18144 36780 18196 36786
rect 18144 36722 18196 36728
rect 18052 36372 18104 36378
rect 18052 36314 18104 36320
rect 17960 36168 18012 36174
rect 17960 36110 18012 36116
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 17776 34944 17828 34950
rect 17776 34886 17828 34892
rect 17684 34060 17736 34066
rect 17684 34002 17736 34008
rect 17590 33552 17646 33561
rect 16948 33516 17000 33522
rect 16948 33458 17000 33464
rect 17408 33516 17460 33522
rect 17590 33487 17646 33496
rect 17408 33458 17460 33464
rect 16856 33380 16908 33386
rect 16856 33322 16908 33328
rect 16868 33114 16896 33322
rect 16856 33108 16908 33114
rect 16856 33050 16908 33056
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 16868 32434 16896 32846
rect 16960 32570 16988 32846
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 17316 32768 17368 32774
rect 17316 32710 17368 32716
rect 16948 32564 17000 32570
rect 16948 32506 17000 32512
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16672 32292 16724 32298
rect 16672 32234 16724 32240
rect 16580 32224 16632 32230
rect 16580 32166 16632 32172
rect 16316 31726 16528 31754
rect 16500 31346 16528 31726
rect 16592 31414 16620 32166
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 16488 31340 16540 31346
rect 16488 31282 16540 31288
rect 16684 31142 16712 32234
rect 16776 31822 16804 32370
rect 16868 31890 16896 32370
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16960 31346 16988 32506
rect 17052 32434 17080 32710
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 17052 32026 17080 32370
rect 17132 32292 17184 32298
rect 17132 32234 17184 32240
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 17144 31906 17172 32234
rect 17328 31906 17356 32710
rect 17420 32570 17448 33458
rect 17500 33448 17552 33454
rect 17500 33390 17552 33396
rect 17512 32978 17540 33390
rect 17500 32972 17552 32978
rect 17500 32914 17552 32920
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17604 32502 17632 33487
rect 17592 32496 17644 32502
rect 17592 32438 17644 32444
rect 17696 32298 17724 34002
rect 17788 33998 17816 34886
rect 17880 34542 17908 35022
rect 17972 34678 18000 36110
rect 18156 35834 18184 36722
rect 18236 36712 18288 36718
rect 18236 36654 18288 36660
rect 18144 35828 18196 35834
rect 18144 35770 18196 35776
rect 18052 35624 18104 35630
rect 18052 35566 18104 35572
rect 17960 34672 18012 34678
rect 17960 34614 18012 34620
rect 17868 34536 17920 34542
rect 17868 34478 17920 34484
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17880 33386 17908 34478
rect 17972 34134 18000 34614
rect 18064 34202 18092 35566
rect 18144 35012 18196 35018
rect 18144 34954 18196 34960
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 17960 34128 18012 34134
rect 17960 34070 18012 34076
rect 18156 34066 18184 34954
rect 18144 34060 18196 34066
rect 18144 34002 18196 34008
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17868 33380 17920 33386
rect 17868 33322 17920 33328
rect 17776 32972 17828 32978
rect 17776 32914 17828 32920
rect 17684 32292 17736 32298
rect 17684 32234 17736 32240
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17052 31878 17172 31906
rect 17236 31878 17356 31906
rect 17512 31906 17540 31962
rect 17684 31952 17736 31958
rect 17512 31878 17632 31906
rect 17684 31894 17736 31900
rect 17052 31482 17080 31878
rect 17236 31770 17264 31878
rect 17144 31742 17264 31770
rect 17316 31816 17368 31822
rect 17316 31758 17368 31764
rect 17500 31816 17552 31822
rect 17500 31758 17552 31764
rect 17040 31476 17092 31482
rect 17040 31418 17092 31424
rect 17144 31346 17172 31742
rect 16948 31340 17000 31346
rect 16948 31282 17000 31288
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 17144 30258 17172 31282
rect 17328 30394 17356 31758
rect 17408 31748 17460 31754
rect 17408 31690 17460 31696
rect 17420 30938 17448 31690
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17512 30734 17540 31758
rect 17500 30728 17552 30734
rect 17500 30670 17552 30676
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 17144 29646 17172 30194
rect 17604 30122 17632 31878
rect 17696 31346 17724 31894
rect 17684 31340 17736 31346
rect 17684 31282 17736 31288
rect 17788 30802 17816 32914
rect 17972 31482 18000 33458
rect 18156 32570 18184 34002
rect 18144 32564 18196 32570
rect 18144 32506 18196 32512
rect 18248 31754 18276 36654
rect 18156 31726 18276 31754
rect 17960 31476 18012 31482
rect 17960 31418 18012 31424
rect 18156 30870 18184 31726
rect 18144 30864 18196 30870
rect 18144 30806 18196 30812
rect 17776 30796 17828 30802
rect 17776 30738 17828 30744
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 17592 30116 17644 30122
rect 17592 30058 17644 30064
rect 17132 29640 17184 29646
rect 17132 29582 17184 29588
rect 16212 28756 16264 28762
rect 16212 28698 16264 28704
rect 15776 27772 16084 27792
rect 15776 27770 15782 27772
rect 15838 27770 15862 27772
rect 15918 27770 15942 27772
rect 15998 27770 16022 27772
rect 16078 27770 16084 27772
rect 15838 27718 15840 27770
rect 16020 27718 16022 27770
rect 15776 27716 15782 27718
rect 15838 27716 15862 27718
rect 15918 27716 15942 27718
rect 15998 27716 16022 27718
rect 16078 27716 16084 27718
rect 15776 27696 16084 27716
rect 15776 26684 16084 26704
rect 15776 26682 15782 26684
rect 15838 26682 15862 26684
rect 15918 26682 15942 26684
rect 15998 26682 16022 26684
rect 16078 26682 16084 26684
rect 15838 26630 15840 26682
rect 16020 26630 16022 26682
rect 15776 26628 15782 26630
rect 15838 26628 15862 26630
rect 15918 26628 15942 26630
rect 15998 26628 16022 26630
rect 16078 26628 16084 26630
rect 15776 26608 16084 26628
rect 15396 26206 15608 26234
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15028 19310 15056 20198
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15396 2650 15424 26206
rect 15776 25596 16084 25616
rect 15776 25594 15782 25596
rect 15838 25594 15862 25596
rect 15918 25594 15942 25596
rect 15998 25594 16022 25596
rect 16078 25594 16084 25596
rect 15838 25542 15840 25594
rect 16020 25542 16022 25594
rect 15776 25540 15782 25542
rect 15838 25540 15862 25542
rect 15918 25540 15942 25542
rect 15998 25540 16022 25542
rect 16078 25540 16084 25542
rect 15776 25520 16084 25540
rect 15776 24508 16084 24528
rect 15776 24506 15782 24508
rect 15838 24506 15862 24508
rect 15918 24506 15942 24508
rect 15998 24506 16022 24508
rect 16078 24506 16084 24508
rect 15838 24454 15840 24506
rect 16020 24454 16022 24506
rect 15776 24452 15782 24454
rect 15838 24452 15862 24454
rect 15918 24452 15942 24454
rect 15998 24452 16022 24454
rect 16078 24452 16084 24454
rect 15776 24432 16084 24452
rect 15776 23420 16084 23440
rect 15776 23418 15782 23420
rect 15838 23418 15862 23420
rect 15918 23418 15942 23420
rect 15998 23418 16022 23420
rect 16078 23418 16084 23420
rect 15838 23366 15840 23418
rect 16020 23366 16022 23418
rect 15776 23364 15782 23366
rect 15838 23364 15862 23366
rect 15918 23364 15942 23366
rect 15998 23364 16022 23366
rect 16078 23364 16084 23366
rect 15776 23344 16084 23364
rect 15776 22332 16084 22352
rect 15776 22330 15782 22332
rect 15838 22330 15862 22332
rect 15918 22330 15942 22332
rect 15998 22330 16022 22332
rect 16078 22330 16084 22332
rect 15838 22278 15840 22330
rect 16020 22278 16022 22330
rect 15776 22276 15782 22278
rect 15838 22276 15862 22278
rect 15918 22276 15942 22278
rect 15998 22276 16022 22278
rect 16078 22276 16084 22278
rect 15776 22256 16084 22276
rect 15776 21244 16084 21264
rect 15776 21242 15782 21244
rect 15838 21242 15862 21244
rect 15918 21242 15942 21244
rect 15998 21242 16022 21244
rect 16078 21242 16084 21244
rect 15838 21190 15840 21242
rect 16020 21190 16022 21242
rect 15776 21188 15782 21190
rect 15838 21188 15862 21190
rect 15918 21188 15942 21190
rect 15998 21188 16022 21190
rect 16078 21188 16084 21190
rect 15776 21168 16084 21188
rect 15776 20156 16084 20176
rect 15776 20154 15782 20156
rect 15838 20154 15862 20156
rect 15918 20154 15942 20156
rect 15998 20154 16022 20156
rect 16078 20154 16084 20156
rect 15838 20102 15840 20154
rect 16020 20102 16022 20154
rect 15776 20100 15782 20102
rect 15838 20100 15862 20102
rect 15918 20100 15942 20102
rect 15998 20100 16022 20102
rect 16078 20100 16084 20102
rect 15776 20080 16084 20100
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15776 19068 16084 19088
rect 15776 19066 15782 19068
rect 15838 19066 15862 19068
rect 15918 19066 15942 19068
rect 15998 19066 16022 19068
rect 16078 19066 16084 19068
rect 15838 19014 15840 19066
rect 16020 19014 16022 19066
rect 15776 19012 15782 19014
rect 15838 19012 15862 19014
rect 15918 19012 15942 19014
rect 15998 19012 16022 19014
rect 16078 19012 16084 19014
rect 15776 18992 16084 19012
rect 15776 17980 16084 18000
rect 15776 17978 15782 17980
rect 15838 17978 15862 17980
rect 15918 17978 15942 17980
rect 15998 17978 16022 17980
rect 16078 17978 16084 17980
rect 15838 17926 15840 17978
rect 16020 17926 16022 17978
rect 15776 17924 15782 17926
rect 15838 17924 15862 17926
rect 15918 17924 15942 17926
rect 15998 17924 16022 17926
rect 16078 17924 16084 17926
rect 15776 17904 16084 17924
rect 15776 16892 16084 16912
rect 15776 16890 15782 16892
rect 15838 16890 15862 16892
rect 15918 16890 15942 16892
rect 15998 16890 16022 16892
rect 16078 16890 16084 16892
rect 15838 16838 15840 16890
rect 16020 16838 16022 16890
rect 15776 16836 15782 16838
rect 15838 16836 15862 16838
rect 15918 16836 15942 16838
rect 15998 16836 16022 16838
rect 16078 16836 16084 16838
rect 15776 16816 16084 16836
rect 15776 15804 16084 15824
rect 15776 15802 15782 15804
rect 15838 15802 15862 15804
rect 15918 15802 15942 15804
rect 15998 15802 16022 15804
rect 16078 15802 16084 15804
rect 15838 15750 15840 15802
rect 16020 15750 16022 15802
rect 15776 15748 15782 15750
rect 15838 15748 15862 15750
rect 15918 15748 15942 15750
rect 15998 15748 16022 15750
rect 16078 15748 16084 15750
rect 15776 15728 16084 15748
rect 15776 14716 16084 14736
rect 15776 14714 15782 14716
rect 15838 14714 15862 14716
rect 15918 14714 15942 14716
rect 15998 14714 16022 14716
rect 16078 14714 16084 14716
rect 15838 14662 15840 14714
rect 16020 14662 16022 14714
rect 15776 14660 15782 14662
rect 15838 14660 15862 14662
rect 15918 14660 15942 14662
rect 15998 14660 16022 14662
rect 16078 14660 16084 14662
rect 15776 14640 16084 14660
rect 15776 13628 16084 13648
rect 15776 13626 15782 13628
rect 15838 13626 15862 13628
rect 15918 13626 15942 13628
rect 15998 13626 16022 13628
rect 16078 13626 16084 13628
rect 15838 13574 15840 13626
rect 16020 13574 16022 13626
rect 15776 13572 15782 13574
rect 15838 13572 15862 13574
rect 15918 13572 15942 13574
rect 15998 13572 16022 13574
rect 16078 13572 16084 13574
rect 15776 13552 16084 13572
rect 15776 12540 16084 12560
rect 15776 12538 15782 12540
rect 15838 12538 15862 12540
rect 15918 12538 15942 12540
rect 15998 12538 16022 12540
rect 16078 12538 16084 12540
rect 15838 12486 15840 12538
rect 16020 12486 16022 12538
rect 15776 12484 15782 12486
rect 15838 12484 15862 12486
rect 15918 12484 15942 12486
rect 15998 12484 16022 12486
rect 16078 12484 16084 12486
rect 15776 12464 16084 12484
rect 15776 11452 16084 11472
rect 15776 11450 15782 11452
rect 15838 11450 15862 11452
rect 15918 11450 15942 11452
rect 15998 11450 16022 11452
rect 16078 11450 16084 11452
rect 15838 11398 15840 11450
rect 16020 11398 16022 11450
rect 15776 11396 15782 11398
rect 15838 11396 15862 11398
rect 15918 11396 15942 11398
rect 15998 11396 16022 11398
rect 16078 11396 16084 11398
rect 15776 11376 16084 11396
rect 15776 10364 16084 10384
rect 15776 10362 15782 10364
rect 15838 10362 15862 10364
rect 15918 10362 15942 10364
rect 15998 10362 16022 10364
rect 16078 10362 16084 10364
rect 15838 10310 15840 10362
rect 16020 10310 16022 10362
rect 15776 10308 15782 10310
rect 15838 10308 15862 10310
rect 15918 10308 15942 10310
rect 15998 10308 16022 10310
rect 16078 10308 16084 10310
rect 15776 10288 16084 10308
rect 15776 9276 16084 9296
rect 15776 9274 15782 9276
rect 15838 9274 15862 9276
rect 15918 9274 15942 9276
rect 15998 9274 16022 9276
rect 16078 9274 16084 9276
rect 15838 9222 15840 9274
rect 16020 9222 16022 9274
rect 15776 9220 15782 9222
rect 15838 9220 15862 9222
rect 15918 9220 15942 9222
rect 15998 9220 16022 9222
rect 16078 9220 16084 9222
rect 15776 9200 16084 9220
rect 15776 8188 16084 8208
rect 15776 8186 15782 8188
rect 15838 8186 15862 8188
rect 15918 8186 15942 8188
rect 15998 8186 16022 8188
rect 16078 8186 16084 8188
rect 15838 8134 15840 8186
rect 16020 8134 16022 8186
rect 15776 8132 15782 8134
rect 15838 8132 15862 8134
rect 15918 8132 15942 8134
rect 15998 8132 16022 8134
rect 16078 8132 16084 8134
rect 15776 8112 16084 8132
rect 15776 7100 16084 7120
rect 15776 7098 15782 7100
rect 15838 7098 15862 7100
rect 15918 7098 15942 7100
rect 15998 7098 16022 7100
rect 16078 7098 16084 7100
rect 15838 7046 15840 7098
rect 16020 7046 16022 7098
rect 15776 7044 15782 7046
rect 15838 7044 15862 7046
rect 15918 7044 15942 7046
rect 15998 7044 16022 7046
rect 16078 7044 16084 7046
rect 15776 7024 16084 7044
rect 15776 6012 16084 6032
rect 15776 6010 15782 6012
rect 15838 6010 15862 6012
rect 15918 6010 15942 6012
rect 15998 6010 16022 6012
rect 16078 6010 16084 6012
rect 15838 5958 15840 6010
rect 16020 5958 16022 6010
rect 15776 5956 15782 5958
rect 15838 5956 15862 5958
rect 15918 5956 15942 5958
rect 15998 5956 16022 5958
rect 16078 5956 16084 5958
rect 15776 5936 16084 5956
rect 15776 4924 16084 4944
rect 15776 4922 15782 4924
rect 15838 4922 15862 4924
rect 15918 4922 15942 4924
rect 15998 4922 16022 4924
rect 16078 4922 16084 4924
rect 15838 4870 15840 4922
rect 16020 4870 16022 4922
rect 15776 4868 15782 4870
rect 15838 4868 15862 4870
rect 15918 4868 15942 4870
rect 15998 4868 16022 4870
rect 16078 4868 16084 4870
rect 15776 4848 16084 4868
rect 15776 3836 16084 3856
rect 15776 3834 15782 3836
rect 15838 3834 15862 3836
rect 15918 3834 15942 3836
rect 15998 3834 16022 3836
rect 16078 3834 16084 3836
rect 15838 3782 15840 3834
rect 16020 3782 16022 3834
rect 15776 3780 15782 3782
rect 15838 3780 15862 3782
rect 15918 3780 15942 3782
rect 15998 3780 16022 3782
rect 16078 3780 16084 3782
rect 15776 3760 16084 3780
rect 16132 3534 16160 19246
rect 17880 16114 17908 30194
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17972 9586 18000 29446
rect 18064 21894 18092 30194
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 18156 28257 18184 28494
rect 18142 28248 18198 28257
rect 18142 28183 18198 28192
rect 18144 22024 18196 22030
rect 18142 21992 18144 22001
rect 18196 21992 18198 22001
rect 18142 21927 18198 21936
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18156 15745 18184 15982
rect 18142 15736 18198 15745
rect 18142 15671 18144 15680
rect 18196 15671 18198 15680
rect 18144 15642 18196 15648
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 18050 9480 18106 9489
rect 18050 9415 18052 9424
rect 18104 9415 18106 9424
rect 18052 9386 18104 9392
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3233 18092 3334
rect 18050 3224 18106 3233
rect 18050 3159 18106 3168
rect 15776 2748 16084 2768
rect 15776 2746 15782 2748
rect 15838 2746 15862 2748
rect 15918 2746 15942 2748
rect 15998 2746 16022 2748
rect 16078 2746 16084 2748
rect 15838 2694 15840 2746
rect 16020 2694 16022 2746
rect 15776 2692 15782 2694
rect 15838 2692 15862 2694
rect 15918 2692 15942 2694
rect 15998 2692 16022 2694
rect 16078 2692 16084 2694
rect 15776 2672 16084 2692
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 12811 2204 13119 2224
rect 12811 2202 12817 2204
rect 12873 2202 12897 2204
rect 12953 2202 12977 2204
rect 13033 2202 13057 2204
rect 13113 2202 13119 2204
rect 12873 2150 12875 2202
rect 13055 2150 13057 2202
rect 12811 2148 12817 2150
rect 12873 2148 12897 2150
rect 12953 2148 12977 2150
rect 13033 2148 13057 2150
rect 13113 2148 13119 2150
rect 12811 2128 13119 2148
rect 17420 800 17448 2382
rect 2502 0 2558 800
rect 7470 0 7526 800
rect 12438 0 12494 800
rect 17406 0 17462 800
<< via2 >>
rect 1490 47252 1546 47288
rect 1490 47232 1492 47252
rect 1492 47232 1544 47252
rect 1544 47232 1546 47252
rect 3921 47354 3977 47356
rect 4001 47354 4057 47356
rect 4081 47354 4137 47356
rect 4161 47354 4217 47356
rect 3921 47302 3967 47354
rect 3967 47302 3977 47354
rect 4001 47302 4031 47354
rect 4031 47302 4043 47354
rect 4043 47302 4057 47354
rect 4081 47302 4095 47354
rect 4095 47302 4107 47354
rect 4107 47302 4137 47354
rect 4161 47302 4171 47354
rect 4171 47302 4217 47354
rect 3921 47300 3977 47302
rect 4001 47300 4057 47302
rect 4081 47300 4137 47302
rect 4161 47300 4217 47302
rect 6886 46810 6942 46812
rect 6966 46810 7022 46812
rect 7046 46810 7102 46812
rect 7126 46810 7182 46812
rect 6886 46758 6932 46810
rect 6932 46758 6942 46810
rect 6966 46758 6996 46810
rect 6996 46758 7008 46810
rect 7008 46758 7022 46810
rect 7046 46758 7060 46810
rect 7060 46758 7072 46810
rect 7072 46758 7102 46810
rect 7126 46758 7136 46810
rect 7136 46758 7182 46810
rect 6886 46756 6942 46758
rect 6966 46756 7022 46758
rect 7046 46756 7102 46758
rect 7126 46756 7182 46758
rect 9852 47354 9908 47356
rect 9932 47354 9988 47356
rect 10012 47354 10068 47356
rect 10092 47354 10148 47356
rect 9852 47302 9898 47354
rect 9898 47302 9908 47354
rect 9932 47302 9962 47354
rect 9962 47302 9974 47354
rect 9974 47302 9988 47354
rect 10012 47302 10026 47354
rect 10026 47302 10038 47354
rect 10038 47302 10068 47354
rect 10092 47302 10102 47354
rect 10102 47302 10148 47354
rect 9852 47300 9908 47302
rect 9932 47300 9988 47302
rect 10012 47300 10068 47302
rect 10092 47300 10148 47302
rect 12817 46810 12873 46812
rect 12897 46810 12953 46812
rect 12977 46810 13033 46812
rect 13057 46810 13113 46812
rect 12817 46758 12863 46810
rect 12863 46758 12873 46810
rect 12897 46758 12927 46810
rect 12927 46758 12939 46810
rect 12939 46758 12953 46810
rect 12977 46758 12991 46810
rect 12991 46758 13003 46810
rect 13003 46758 13033 46810
rect 13057 46758 13067 46810
rect 13067 46758 13113 46810
rect 12817 46756 12873 46758
rect 12897 46756 12953 46758
rect 12977 46756 13033 46758
rect 13057 46756 13113 46758
rect 3921 46266 3977 46268
rect 4001 46266 4057 46268
rect 4081 46266 4137 46268
rect 4161 46266 4217 46268
rect 3921 46214 3967 46266
rect 3967 46214 3977 46266
rect 4001 46214 4031 46266
rect 4031 46214 4043 46266
rect 4043 46214 4057 46266
rect 4081 46214 4095 46266
rect 4095 46214 4107 46266
rect 4107 46214 4137 46266
rect 4161 46214 4171 46266
rect 4171 46214 4217 46266
rect 3921 46212 3977 46214
rect 4001 46212 4057 46214
rect 4081 46212 4137 46214
rect 4161 46212 4217 46214
rect 9852 46266 9908 46268
rect 9932 46266 9988 46268
rect 10012 46266 10068 46268
rect 10092 46266 10148 46268
rect 9852 46214 9898 46266
rect 9898 46214 9908 46266
rect 9932 46214 9962 46266
rect 9962 46214 9974 46266
rect 9974 46214 9988 46266
rect 10012 46214 10026 46266
rect 10026 46214 10038 46266
rect 10038 46214 10068 46266
rect 10092 46214 10102 46266
rect 10102 46214 10148 46266
rect 9852 46212 9908 46214
rect 9932 46212 9988 46214
rect 10012 46212 10068 46214
rect 10092 46212 10148 46214
rect 1490 41656 1546 41712
rect 1858 36100 1914 36136
rect 1858 36080 1860 36100
rect 1860 36080 1912 36100
rect 1912 36080 1914 36100
rect 6886 45722 6942 45724
rect 6966 45722 7022 45724
rect 7046 45722 7102 45724
rect 7126 45722 7182 45724
rect 6886 45670 6932 45722
rect 6932 45670 6942 45722
rect 6966 45670 6996 45722
rect 6996 45670 7008 45722
rect 7008 45670 7022 45722
rect 7046 45670 7060 45722
rect 7060 45670 7072 45722
rect 7072 45670 7102 45722
rect 7126 45670 7136 45722
rect 7136 45670 7182 45722
rect 6886 45668 6942 45670
rect 6966 45668 7022 45670
rect 7046 45668 7102 45670
rect 7126 45668 7182 45670
rect 12817 45722 12873 45724
rect 12897 45722 12953 45724
rect 12977 45722 13033 45724
rect 13057 45722 13113 45724
rect 12817 45670 12863 45722
rect 12863 45670 12873 45722
rect 12897 45670 12927 45722
rect 12927 45670 12939 45722
rect 12939 45670 12953 45722
rect 12977 45670 12991 45722
rect 12991 45670 13003 45722
rect 13003 45670 13033 45722
rect 13057 45670 13067 45722
rect 13067 45670 13113 45722
rect 12817 45668 12873 45670
rect 12897 45668 12953 45670
rect 12977 45668 13033 45670
rect 13057 45668 13113 45670
rect 3921 45178 3977 45180
rect 4001 45178 4057 45180
rect 4081 45178 4137 45180
rect 4161 45178 4217 45180
rect 3921 45126 3967 45178
rect 3967 45126 3977 45178
rect 4001 45126 4031 45178
rect 4031 45126 4043 45178
rect 4043 45126 4057 45178
rect 4081 45126 4095 45178
rect 4095 45126 4107 45178
rect 4107 45126 4137 45178
rect 4161 45126 4171 45178
rect 4171 45126 4217 45178
rect 3921 45124 3977 45126
rect 4001 45124 4057 45126
rect 4081 45124 4137 45126
rect 4161 45124 4217 45126
rect 9852 45178 9908 45180
rect 9932 45178 9988 45180
rect 10012 45178 10068 45180
rect 10092 45178 10148 45180
rect 9852 45126 9898 45178
rect 9898 45126 9908 45178
rect 9932 45126 9962 45178
rect 9962 45126 9974 45178
rect 9974 45126 9988 45178
rect 10012 45126 10026 45178
rect 10026 45126 10038 45178
rect 10038 45126 10068 45178
rect 10092 45126 10102 45178
rect 10102 45126 10148 45178
rect 9852 45124 9908 45126
rect 9932 45124 9988 45126
rect 10012 45124 10068 45126
rect 10092 45124 10148 45126
rect 6886 44634 6942 44636
rect 6966 44634 7022 44636
rect 7046 44634 7102 44636
rect 7126 44634 7182 44636
rect 6886 44582 6932 44634
rect 6932 44582 6942 44634
rect 6966 44582 6996 44634
rect 6996 44582 7008 44634
rect 7008 44582 7022 44634
rect 7046 44582 7060 44634
rect 7060 44582 7072 44634
rect 7072 44582 7102 44634
rect 7126 44582 7136 44634
rect 7136 44582 7182 44634
rect 6886 44580 6942 44582
rect 6966 44580 7022 44582
rect 7046 44580 7102 44582
rect 7126 44580 7182 44582
rect 12817 44634 12873 44636
rect 12897 44634 12953 44636
rect 12977 44634 13033 44636
rect 13057 44634 13113 44636
rect 12817 44582 12863 44634
rect 12863 44582 12873 44634
rect 12897 44582 12927 44634
rect 12927 44582 12939 44634
rect 12939 44582 12953 44634
rect 12977 44582 12991 44634
rect 12991 44582 13003 44634
rect 13003 44582 13033 44634
rect 13057 44582 13067 44634
rect 13067 44582 13113 44634
rect 12817 44580 12873 44582
rect 12897 44580 12953 44582
rect 12977 44580 13033 44582
rect 13057 44580 13113 44582
rect 3921 44090 3977 44092
rect 4001 44090 4057 44092
rect 4081 44090 4137 44092
rect 4161 44090 4217 44092
rect 3921 44038 3967 44090
rect 3967 44038 3977 44090
rect 4001 44038 4031 44090
rect 4031 44038 4043 44090
rect 4043 44038 4057 44090
rect 4081 44038 4095 44090
rect 4095 44038 4107 44090
rect 4107 44038 4137 44090
rect 4161 44038 4171 44090
rect 4171 44038 4217 44090
rect 3921 44036 3977 44038
rect 4001 44036 4057 44038
rect 4081 44036 4137 44038
rect 4161 44036 4217 44038
rect 9852 44090 9908 44092
rect 9932 44090 9988 44092
rect 10012 44090 10068 44092
rect 10092 44090 10148 44092
rect 9852 44038 9898 44090
rect 9898 44038 9908 44090
rect 9932 44038 9962 44090
rect 9962 44038 9974 44090
rect 9974 44038 9988 44090
rect 10012 44038 10026 44090
rect 10026 44038 10038 44090
rect 10038 44038 10068 44090
rect 10092 44038 10102 44090
rect 10102 44038 10148 44090
rect 9852 44036 9908 44038
rect 9932 44036 9988 44038
rect 10012 44036 10068 44038
rect 10092 44036 10148 44038
rect 6886 43546 6942 43548
rect 6966 43546 7022 43548
rect 7046 43546 7102 43548
rect 7126 43546 7182 43548
rect 6886 43494 6932 43546
rect 6932 43494 6942 43546
rect 6966 43494 6996 43546
rect 6996 43494 7008 43546
rect 7008 43494 7022 43546
rect 7046 43494 7060 43546
rect 7060 43494 7072 43546
rect 7072 43494 7102 43546
rect 7126 43494 7136 43546
rect 7136 43494 7182 43546
rect 6886 43492 6942 43494
rect 6966 43492 7022 43494
rect 7046 43492 7102 43494
rect 7126 43492 7182 43494
rect 12817 43546 12873 43548
rect 12897 43546 12953 43548
rect 12977 43546 13033 43548
rect 13057 43546 13113 43548
rect 12817 43494 12863 43546
rect 12863 43494 12873 43546
rect 12897 43494 12927 43546
rect 12927 43494 12939 43546
rect 12939 43494 12953 43546
rect 12977 43494 12991 43546
rect 12991 43494 13003 43546
rect 13003 43494 13033 43546
rect 13057 43494 13067 43546
rect 13067 43494 13113 43546
rect 12817 43492 12873 43494
rect 12897 43492 12953 43494
rect 12977 43492 13033 43494
rect 13057 43492 13113 43494
rect 3921 43002 3977 43004
rect 4001 43002 4057 43004
rect 4081 43002 4137 43004
rect 4161 43002 4217 43004
rect 3921 42950 3967 43002
rect 3967 42950 3977 43002
rect 4001 42950 4031 43002
rect 4031 42950 4043 43002
rect 4043 42950 4057 43002
rect 4081 42950 4095 43002
rect 4095 42950 4107 43002
rect 4107 42950 4137 43002
rect 4161 42950 4171 43002
rect 4171 42950 4217 43002
rect 3921 42948 3977 42950
rect 4001 42948 4057 42950
rect 4081 42948 4137 42950
rect 4161 42948 4217 42950
rect 9852 43002 9908 43004
rect 9932 43002 9988 43004
rect 10012 43002 10068 43004
rect 10092 43002 10148 43004
rect 9852 42950 9898 43002
rect 9898 42950 9908 43002
rect 9932 42950 9962 43002
rect 9962 42950 9974 43002
rect 9974 42950 9988 43002
rect 10012 42950 10026 43002
rect 10026 42950 10038 43002
rect 10038 42950 10068 43002
rect 10092 42950 10102 43002
rect 10102 42950 10148 43002
rect 9852 42948 9908 42950
rect 9932 42948 9988 42950
rect 10012 42948 10068 42950
rect 10092 42948 10148 42950
rect 6886 42458 6942 42460
rect 6966 42458 7022 42460
rect 7046 42458 7102 42460
rect 7126 42458 7182 42460
rect 6886 42406 6932 42458
rect 6932 42406 6942 42458
rect 6966 42406 6996 42458
rect 6996 42406 7008 42458
rect 7008 42406 7022 42458
rect 7046 42406 7060 42458
rect 7060 42406 7072 42458
rect 7072 42406 7102 42458
rect 7126 42406 7136 42458
rect 7136 42406 7182 42458
rect 6886 42404 6942 42406
rect 6966 42404 7022 42406
rect 7046 42404 7102 42406
rect 7126 42404 7182 42406
rect 12817 42458 12873 42460
rect 12897 42458 12953 42460
rect 12977 42458 13033 42460
rect 13057 42458 13113 42460
rect 12817 42406 12863 42458
rect 12863 42406 12873 42458
rect 12897 42406 12927 42458
rect 12927 42406 12939 42458
rect 12939 42406 12953 42458
rect 12977 42406 12991 42458
rect 12991 42406 13003 42458
rect 13003 42406 13033 42458
rect 13057 42406 13067 42458
rect 13067 42406 13113 42458
rect 12817 42404 12873 42406
rect 12897 42404 12953 42406
rect 12977 42404 13033 42406
rect 13057 42404 13113 42406
rect 3921 41914 3977 41916
rect 4001 41914 4057 41916
rect 4081 41914 4137 41916
rect 4161 41914 4217 41916
rect 3921 41862 3967 41914
rect 3967 41862 3977 41914
rect 4001 41862 4031 41914
rect 4031 41862 4043 41914
rect 4043 41862 4057 41914
rect 4081 41862 4095 41914
rect 4095 41862 4107 41914
rect 4107 41862 4137 41914
rect 4161 41862 4171 41914
rect 4171 41862 4217 41914
rect 3921 41860 3977 41862
rect 4001 41860 4057 41862
rect 4081 41860 4137 41862
rect 4161 41860 4217 41862
rect 9852 41914 9908 41916
rect 9932 41914 9988 41916
rect 10012 41914 10068 41916
rect 10092 41914 10148 41916
rect 9852 41862 9898 41914
rect 9898 41862 9908 41914
rect 9932 41862 9962 41914
rect 9962 41862 9974 41914
rect 9974 41862 9988 41914
rect 10012 41862 10026 41914
rect 10026 41862 10038 41914
rect 10038 41862 10068 41914
rect 10092 41862 10102 41914
rect 10102 41862 10148 41914
rect 9852 41860 9908 41862
rect 9932 41860 9988 41862
rect 10012 41860 10068 41862
rect 10092 41860 10148 41862
rect 6886 41370 6942 41372
rect 6966 41370 7022 41372
rect 7046 41370 7102 41372
rect 7126 41370 7182 41372
rect 6886 41318 6932 41370
rect 6932 41318 6942 41370
rect 6966 41318 6996 41370
rect 6996 41318 7008 41370
rect 7008 41318 7022 41370
rect 7046 41318 7060 41370
rect 7060 41318 7072 41370
rect 7072 41318 7102 41370
rect 7126 41318 7136 41370
rect 7136 41318 7182 41370
rect 6886 41316 6942 41318
rect 6966 41316 7022 41318
rect 7046 41316 7102 41318
rect 7126 41316 7182 41318
rect 12817 41370 12873 41372
rect 12897 41370 12953 41372
rect 12977 41370 13033 41372
rect 13057 41370 13113 41372
rect 12817 41318 12863 41370
rect 12863 41318 12873 41370
rect 12897 41318 12927 41370
rect 12927 41318 12939 41370
rect 12939 41318 12953 41370
rect 12977 41318 12991 41370
rect 12991 41318 13003 41370
rect 13003 41318 13033 41370
rect 13057 41318 13067 41370
rect 13067 41318 13113 41370
rect 12817 41316 12873 41318
rect 12897 41316 12953 41318
rect 12977 41316 13033 41318
rect 13057 41316 13113 41318
rect 3921 40826 3977 40828
rect 4001 40826 4057 40828
rect 4081 40826 4137 40828
rect 4161 40826 4217 40828
rect 3921 40774 3967 40826
rect 3967 40774 3977 40826
rect 4001 40774 4031 40826
rect 4031 40774 4043 40826
rect 4043 40774 4057 40826
rect 4081 40774 4095 40826
rect 4095 40774 4107 40826
rect 4107 40774 4137 40826
rect 4161 40774 4171 40826
rect 4171 40774 4217 40826
rect 3921 40772 3977 40774
rect 4001 40772 4057 40774
rect 4081 40772 4137 40774
rect 4161 40772 4217 40774
rect 9852 40826 9908 40828
rect 9932 40826 9988 40828
rect 10012 40826 10068 40828
rect 10092 40826 10148 40828
rect 9852 40774 9898 40826
rect 9898 40774 9908 40826
rect 9932 40774 9962 40826
rect 9962 40774 9974 40826
rect 9974 40774 9988 40826
rect 10012 40774 10026 40826
rect 10026 40774 10038 40826
rect 10038 40774 10068 40826
rect 10092 40774 10102 40826
rect 10102 40774 10148 40826
rect 9852 40772 9908 40774
rect 9932 40772 9988 40774
rect 10012 40772 10068 40774
rect 10092 40772 10148 40774
rect 6886 40282 6942 40284
rect 6966 40282 7022 40284
rect 7046 40282 7102 40284
rect 7126 40282 7182 40284
rect 6886 40230 6932 40282
rect 6932 40230 6942 40282
rect 6966 40230 6996 40282
rect 6996 40230 7008 40282
rect 7008 40230 7022 40282
rect 7046 40230 7060 40282
rect 7060 40230 7072 40282
rect 7072 40230 7102 40282
rect 7126 40230 7136 40282
rect 7136 40230 7182 40282
rect 6886 40228 6942 40230
rect 6966 40228 7022 40230
rect 7046 40228 7102 40230
rect 7126 40228 7182 40230
rect 12817 40282 12873 40284
rect 12897 40282 12953 40284
rect 12977 40282 13033 40284
rect 13057 40282 13113 40284
rect 12817 40230 12863 40282
rect 12863 40230 12873 40282
rect 12897 40230 12927 40282
rect 12927 40230 12939 40282
rect 12939 40230 12953 40282
rect 12977 40230 12991 40282
rect 12991 40230 13003 40282
rect 13003 40230 13033 40282
rect 13057 40230 13067 40282
rect 13067 40230 13113 40282
rect 12817 40228 12873 40230
rect 12897 40228 12953 40230
rect 12977 40228 13033 40230
rect 13057 40228 13113 40230
rect 3921 39738 3977 39740
rect 4001 39738 4057 39740
rect 4081 39738 4137 39740
rect 4161 39738 4217 39740
rect 3921 39686 3967 39738
rect 3967 39686 3977 39738
rect 4001 39686 4031 39738
rect 4031 39686 4043 39738
rect 4043 39686 4057 39738
rect 4081 39686 4095 39738
rect 4095 39686 4107 39738
rect 4107 39686 4137 39738
rect 4161 39686 4171 39738
rect 4171 39686 4217 39738
rect 3921 39684 3977 39686
rect 4001 39684 4057 39686
rect 4081 39684 4137 39686
rect 4161 39684 4217 39686
rect 9852 39738 9908 39740
rect 9932 39738 9988 39740
rect 10012 39738 10068 39740
rect 10092 39738 10148 39740
rect 9852 39686 9898 39738
rect 9898 39686 9908 39738
rect 9932 39686 9962 39738
rect 9962 39686 9974 39738
rect 9974 39686 9988 39738
rect 10012 39686 10026 39738
rect 10026 39686 10038 39738
rect 10038 39686 10068 39738
rect 10092 39686 10102 39738
rect 10102 39686 10148 39738
rect 9852 39684 9908 39686
rect 9932 39684 9988 39686
rect 10012 39684 10068 39686
rect 10092 39684 10148 39686
rect 6886 39194 6942 39196
rect 6966 39194 7022 39196
rect 7046 39194 7102 39196
rect 7126 39194 7182 39196
rect 6886 39142 6932 39194
rect 6932 39142 6942 39194
rect 6966 39142 6996 39194
rect 6996 39142 7008 39194
rect 7008 39142 7022 39194
rect 7046 39142 7060 39194
rect 7060 39142 7072 39194
rect 7072 39142 7102 39194
rect 7126 39142 7136 39194
rect 7136 39142 7182 39194
rect 6886 39140 6942 39142
rect 6966 39140 7022 39142
rect 7046 39140 7102 39142
rect 7126 39140 7182 39142
rect 12817 39194 12873 39196
rect 12897 39194 12953 39196
rect 12977 39194 13033 39196
rect 13057 39194 13113 39196
rect 12817 39142 12863 39194
rect 12863 39142 12873 39194
rect 12897 39142 12927 39194
rect 12927 39142 12939 39194
rect 12939 39142 12953 39194
rect 12977 39142 12991 39194
rect 12991 39142 13003 39194
rect 13003 39142 13033 39194
rect 13057 39142 13067 39194
rect 13067 39142 13113 39194
rect 12817 39140 12873 39142
rect 12897 39140 12953 39142
rect 12977 39140 13033 39142
rect 13057 39140 13113 39142
rect 3921 38650 3977 38652
rect 4001 38650 4057 38652
rect 4081 38650 4137 38652
rect 4161 38650 4217 38652
rect 3921 38598 3967 38650
rect 3967 38598 3977 38650
rect 4001 38598 4031 38650
rect 4031 38598 4043 38650
rect 4043 38598 4057 38650
rect 4081 38598 4095 38650
rect 4095 38598 4107 38650
rect 4107 38598 4137 38650
rect 4161 38598 4171 38650
rect 4171 38598 4217 38650
rect 3921 38596 3977 38598
rect 4001 38596 4057 38598
rect 4081 38596 4137 38598
rect 4161 38596 4217 38598
rect 9852 38650 9908 38652
rect 9932 38650 9988 38652
rect 10012 38650 10068 38652
rect 10092 38650 10148 38652
rect 9852 38598 9898 38650
rect 9898 38598 9908 38650
rect 9932 38598 9962 38650
rect 9962 38598 9974 38650
rect 9974 38598 9988 38650
rect 10012 38598 10026 38650
rect 10026 38598 10038 38650
rect 10038 38598 10068 38650
rect 10092 38598 10102 38650
rect 10102 38598 10148 38650
rect 9852 38596 9908 38598
rect 9932 38596 9988 38598
rect 10012 38596 10068 38598
rect 10092 38596 10148 38598
rect 6886 38106 6942 38108
rect 6966 38106 7022 38108
rect 7046 38106 7102 38108
rect 7126 38106 7182 38108
rect 6886 38054 6932 38106
rect 6932 38054 6942 38106
rect 6966 38054 6996 38106
rect 6996 38054 7008 38106
rect 7008 38054 7022 38106
rect 7046 38054 7060 38106
rect 7060 38054 7072 38106
rect 7072 38054 7102 38106
rect 7126 38054 7136 38106
rect 7136 38054 7182 38106
rect 6886 38052 6942 38054
rect 6966 38052 7022 38054
rect 7046 38052 7102 38054
rect 7126 38052 7182 38054
rect 12817 38106 12873 38108
rect 12897 38106 12953 38108
rect 12977 38106 13033 38108
rect 13057 38106 13113 38108
rect 12817 38054 12863 38106
rect 12863 38054 12873 38106
rect 12897 38054 12927 38106
rect 12927 38054 12939 38106
rect 12939 38054 12953 38106
rect 12977 38054 12991 38106
rect 12991 38054 13003 38106
rect 13003 38054 13033 38106
rect 13057 38054 13067 38106
rect 13067 38054 13113 38106
rect 12817 38052 12873 38054
rect 12897 38052 12953 38054
rect 12977 38052 13033 38054
rect 13057 38052 13113 38054
rect 3921 37562 3977 37564
rect 4001 37562 4057 37564
rect 4081 37562 4137 37564
rect 4161 37562 4217 37564
rect 3921 37510 3967 37562
rect 3967 37510 3977 37562
rect 4001 37510 4031 37562
rect 4031 37510 4043 37562
rect 4043 37510 4057 37562
rect 4081 37510 4095 37562
rect 4095 37510 4107 37562
rect 4107 37510 4137 37562
rect 4161 37510 4171 37562
rect 4171 37510 4217 37562
rect 3921 37508 3977 37510
rect 4001 37508 4057 37510
rect 4081 37508 4137 37510
rect 4161 37508 4217 37510
rect 9852 37562 9908 37564
rect 9932 37562 9988 37564
rect 10012 37562 10068 37564
rect 10092 37562 10148 37564
rect 9852 37510 9898 37562
rect 9898 37510 9908 37562
rect 9932 37510 9962 37562
rect 9962 37510 9974 37562
rect 9974 37510 9988 37562
rect 10012 37510 10026 37562
rect 10026 37510 10038 37562
rect 10038 37510 10068 37562
rect 10092 37510 10102 37562
rect 10102 37510 10148 37562
rect 9852 37508 9908 37510
rect 9932 37508 9988 37510
rect 10012 37508 10068 37510
rect 10092 37508 10148 37510
rect 6886 37018 6942 37020
rect 6966 37018 7022 37020
rect 7046 37018 7102 37020
rect 7126 37018 7182 37020
rect 6886 36966 6932 37018
rect 6932 36966 6942 37018
rect 6966 36966 6996 37018
rect 6996 36966 7008 37018
rect 7008 36966 7022 37018
rect 7046 36966 7060 37018
rect 7060 36966 7072 37018
rect 7072 36966 7102 37018
rect 7126 36966 7136 37018
rect 7136 36966 7182 37018
rect 6886 36964 6942 36966
rect 6966 36964 7022 36966
rect 7046 36964 7102 36966
rect 7126 36964 7182 36966
rect 12817 37018 12873 37020
rect 12897 37018 12953 37020
rect 12977 37018 13033 37020
rect 13057 37018 13113 37020
rect 12817 36966 12863 37018
rect 12863 36966 12873 37018
rect 12897 36966 12927 37018
rect 12927 36966 12939 37018
rect 12939 36966 12953 37018
rect 12977 36966 12991 37018
rect 12991 36966 13003 37018
rect 13003 36966 13033 37018
rect 13057 36966 13067 37018
rect 13067 36966 13113 37018
rect 12817 36964 12873 36966
rect 12897 36964 12953 36966
rect 12977 36964 13033 36966
rect 13057 36964 13113 36966
rect 3921 36474 3977 36476
rect 4001 36474 4057 36476
rect 4081 36474 4137 36476
rect 4161 36474 4217 36476
rect 3921 36422 3967 36474
rect 3967 36422 3977 36474
rect 4001 36422 4031 36474
rect 4031 36422 4043 36474
rect 4043 36422 4057 36474
rect 4081 36422 4095 36474
rect 4095 36422 4107 36474
rect 4107 36422 4137 36474
rect 4161 36422 4171 36474
rect 4171 36422 4217 36474
rect 3921 36420 3977 36422
rect 4001 36420 4057 36422
rect 4081 36420 4137 36422
rect 4161 36420 4217 36422
rect 9852 36474 9908 36476
rect 9932 36474 9988 36476
rect 10012 36474 10068 36476
rect 10092 36474 10148 36476
rect 9852 36422 9898 36474
rect 9898 36422 9908 36474
rect 9932 36422 9962 36474
rect 9962 36422 9974 36474
rect 9974 36422 9988 36474
rect 10012 36422 10026 36474
rect 10026 36422 10038 36474
rect 10038 36422 10068 36474
rect 10092 36422 10102 36474
rect 10102 36422 10148 36474
rect 9852 36420 9908 36422
rect 9932 36420 9988 36422
rect 10012 36420 10068 36422
rect 10092 36420 10148 36422
rect 6886 35930 6942 35932
rect 6966 35930 7022 35932
rect 7046 35930 7102 35932
rect 7126 35930 7182 35932
rect 6886 35878 6932 35930
rect 6932 35878 6942 35930
rect 6966 35878 6996 35930
rect 6996 35878 7008 35930
rect 7008 35878 7022 35930
rect 7046 35878 7060 35930
rect 7060 35878 7072 35930
rect 7072 35878 7102 35930
rect 7126 35878 7136 35930
rect 7136 35878 7182 35930
rect 6886 35876 6942 35878
rect 6966 35876 7022 35878
rect 7046 35876 7102 35878
rect 7126 35876 7182 35878
rect 12817 35930 12873 35932
rect 12897 35930 12953 35932
rect 12977 35930 13033 35932
rect 13057 35930 13113 35932
rect 12817 35878 12863 35930
rect 12863 35878 12873 35930
rect 12897 35878 12927 35930
rect 12927 35878 12939 35930
rect 12939 35878 12953 35930
rect 12977 35878 12991 35930
rect 12991 35878 13003 35930
rect 13003 35878 13033 35930
rect 13057 35878 13067 35930
rect 13067 35878 13113 35930
rect 12817 35876 12873 35878
rect 12897 35876 12953 35878
rect 12977 35876 13033 35878
rect 13057 35876 13113 35878
rect 3921 35386 3977 35388
rect 4001 35386 4057 35388
rect 4081 35386 4137 35388
rect 4161 35386 4217 35388
rect 3921 35334 3967 35386
rect 3967 35334 3977 35386
rect 4001 35334 4031 35386
rect 4031 35334 4043 35386
rect 4043 35334 4057 35386
rect 4081 35334 4095 35386
rect 4095 35334 4107 35386
rect 4107 35334 4137 35386
rect 4161 35334 4171 35386
rect 4171 35334 4217 35386
rect 3921 35332 3977 35334
rect 4001 35332 4057 35334
rect 4081 35332 4137 35334
rect 4161 35332 4217 35334
rect 9852 35386 9908 35388
rect 9932 35386 9988 35388
rect 10012 35386 10068 35388
rect 10092 35386 10148 35388
rect 9852 35334 9898 35386
rect 9898 35334 9908 35386
rect 9932 35334 9962 35386
rect 9962 35334 9974 35386
rect 9974 35334 9988 35386
rect 10012 35334 10026 35386
rect 10026 35334 10038 35386
rect 10038 35334 10068 35386
rect 10092 35334 10102 35386
rect 10102 35334 10148 35386
rect 9852 35332 9908 35334
rect 9932 35332 9988 35334
rect 10012 35332 10068 35334
rect 10092 35332 10148 35334
rect 6886 34842 6942 34844
rect 6966 34842 7022 34844
rect 7046 34842 7102 34844
rect 7126 34842 7182 34844
rect 6886 34790 6932 34842
rect 6932 34790 6942 34842
rect 6966 34790 6996 34842
rect 6996 34790 7008 34842
rect 7008 34790 7022 34842
rect 7046 34790 7060 34842
rect 7060 34790 7072 34842
rect 7072 34790 7102 34842
rect 7126 34790 7136 34842
rect 7136 34790 7182 34842
rect 6886 34788 6942 34790
rect 6966 34788 7022 34790
rect 7046 34788 7102 34790
rect 7126 34788 7182 34790
rect 12817 34842 12873 34844
rect 12897 34842 12953 34844
rect 12977 34842 13033 34844
rect 13057 34842 13113 34844
rect 12817 34790 12863 34842
rect 12863 34790 12873 34842
rect 12897 34790 12927 34842
rect 12927 34790 12939 34842
rect 12939 34790 12953 34842
rect 12977 34790 12991 34842
rect 12991 34790 13003 34842
rect 13003 34790 13033 34842
rect 13057 34790 13067 34842
rect 13067 34790 13113 34842
rect 12817 34788 12873 34790
rect 12897 34788 12953 34790
rect 12977 34788 13033 34790
rect 13057 34788 13113 34790
rect 3921 34298 3977 34300
rect 4001 34298 4057 34300
rect 4081 34298 4137 34300
rect 4161 34298 4217 34300
rect 3921 34246 3967 34298
rect 3967 34246 3977 34298
rect 4001 34246 4031 34298
rect 4031 34246 4043 34298
rect 4043 34246 4057 34298
rect 4081 34246 4095 34298
rect 4095 34246 4107 34298
rect 4107 34246 4137 34298
rect 4161 34246 4171 34298
rect 4171 34246 4217 34298
rect 3921 34244 3977 34246
rect 4001 34244 4057 34246
rect 4081 34244 4137 34246
rect 4161 34244 4217 34246
rect 9852 34298 9908 34300
rect 9932 34298 9988 34300
rect 10012 34298 10068 34300
rect 10092 34298 10148 34300
rect 9852 34246 9898 34298
rect 9898 34246 9908 34298
rect 9932 34246 9962 34298
rect 9962 34246 9974 34298
rect 9974 34246 9988 34298
rect 10012 34246 10026 34298
rect 10026 34246 10038 34298
rect 10038 34246 10068 34298
rect 10092 34246 10102 34298
rect 10102 34246 10148 34298
rect 9852 34244 9908 34246
rect 9932 34244 9988 34246
rect 10012 34244 10068 34246
rect 10092 34244 10148 34246
rect 6886 33754 6942 33756
rect 6966 33754 7022 33756
rect 7046 33754 7102 33756
rect 7126 33754 7182 33756
rect 6886 33702 6932 33754
rect 6932 33702 6942 33754
rect 6966 33702 6996 33754
rect 6996 33702 7008 33754
rect 7008 33702 7022 33754
rect 7046 33702 7060 33754
rect 7060 33702 7072 33754
rect 7072 33702 7102 33754
rect 7126 33702 7136 33754
rect 7136 33702 7182 33754
rect 6886 33700 6942 33702
rect 6966 33700 7022 33702
rect 7046 33700 7102 33702
rect 7126 33700 7182 33702
rect 3921 33210 3977 33212
rect 4001 33210 4057 33212
rect 4081 33210 4137 33212
rect 4161 33210 4217 33212
rect 3921 33158 3967 33210
rect 3967 33158 3977 33210
rect 4001 33158 4031 33210
rect 4031 33158 4043 33210
rect 4043 33158 4057 33210
rect 4081 33158 4095 33210
rect 4095 33158 4107 33210
rect 4107 33158 4137 33210
rect 4161 33158 4171 33210
rect 4171 33158 4217 33210
rect 3921 33156 3977 33158
rect 4001 33156 4057 33158
rect 4081 33156 4137 33158
rect 4161 33156 4217 33158
rect 9852 33210 9908 33212
rect 9932 33210 9988 33212
rect 10012 33210 10068 33212
rect 10092 33210 10148 33212
rect 9852 33158 9898 33210
rect 9898 33158 9908 33210
rect 9932 33158 9962 33210
rect 9962 33158 9974 33210
rect 9974 33158 9988 33210
rect 10012 33158 10026 33210
rect 10026 33158 10038 33210
rect 10038 33158 10068 33210
rect 10092 33158 10102 33210
rect 10102 33158 10148 33210
rect 9852 33156 9908 33158
rect 9932 33156 9988 33158
rect 10012 33156 10068 33158
rect 10092 33156 10148 33158
rect 12817 33754 12873 33756
rect 12897 33754 12953 33756
rect 12977 33754 13033 33756
rect 13057 33754 13113 33756
rect 12817 33702 12863 33754
rect 12863 33702 12873 33754
rect 12897 33702 12927 33754
rect 12927 33702 12939 33754
rect 12939 33702 12953 33754
rect 12977 33702 12991 33754
rect 12991 33702 13003 33754
rect 13003 33702 13033 33754
rect 13057 33702 13067 33754
rect 13067 33702 13113 33754
rect 12817 33700 12873 33702
rect 12897 33700 12953 33702
rect 12977 33700 13033 33702
rect 13057 33700 13113 33702
rect 13542 33516 13598 33552
rect 13542 33496 13544 33516
rect 13544 33496 13596 33516
rect 13596 33496 13598 33516
rect 6886 32666 6942 32668
rect 6966 32666 7022 32668
rect 7046 32666 7102 32668
rect 7126 32666 7182 32668
rect 6886 32614 6932 32666
rect 6932 32614 6942 32666
rect 6966 32614 6996 32666
rect 6996 32614 7008 32666
rect 7008 32614 7022 32666
rect 7046 32614 7060 32666
rect 7060 32614 7072 32666
rect 7072 32614 7102 32666
rect 7126 32614 7136 32666
rect 7136 32614 7182 32666
rect 6886 32612 6942 32614
rect 6966 32612 7022 32614
rect 7046 32612 7102 32614
rect 7126 32612 7182 32614
rect 3921 32122 3977 32124
rect 4001 32122 4057 32124
rect 4081 32122 4137 32124
rect 4161 32122 4217 32124
rect 3921 32070 3967 32122
rect 3967 32070 3977 32122
rect 4001 32070 4031 32122
rect 4031 32070 4043 32122
rect 4043 32070 4057 32122
rect 4081 32070 4095 32122
rect 4095 32070 4107 32122
rect 4107 32070 4137 32122
rect 4161 32070 4171 32122
rect 4171 32070 4217 32122
rect 3921 32068 3977 32070
rect 4001 32068 4057 32070
rect 4081 32068 4137 32070
rect 4161 32068 4217 32070
rect 9852 32122 9908 32124
rect 9932 32122 9988 32124
rect 10012 32122 10068 32124
rect 10092 32122 10148 32124
rect 9852 32070 9898 32122
rect 9898 32070 9908 32122
rect 9932 32070 9962 32122
rect 9962 32070 9974 32122
rect 9974 32070 9988 32122
rect 10012 32070 10026 32122
rect 10026 32070 10038 32122
rect 10038 32070 10068 32122
rect 10092 32070 10102 32122
rect 10102 32070 10148 32122
rect 9852 32068 9908 32070
rect 9932 32068 9988 32070
rect 10012 32068 10068 32070
rect 10092 32068 10148 32070
rect 6886 31578 6942 31580
rect 6966 31578 7022 31580
rect 7046 31578 7102 31580
rect 7126 31578 7182 31580
rect 6886 31526 6932 31578
rect 6932 31526 6942 31578
rect 6966 31526 6996 31578
rect 6996 31526 7008 31578
rect 7008 31526 7022 31578
rect 7046 31526 7060 31578
rect 7060 31526 7072 31578
rect 7072 31526 7102 31578
rect 7126 31526 7136 31578
rect 7136 31526 7182 31578
rect 6886 31524 6942 31526
rect 6966 31524 7022 31526
rect 7046 31524 7102 31526
rect 7126 31524 7182 31526
rect 12817 32666 12873 32668
rect 12897 32666 12953 32668
rect 12977 32666 13033 32668
rect 13057 32666 13113 32668
rect 12817 32614 12863 32666
rect 12863 32614 12873 32666
rect 12897 32614 12927 32666
rect 12927 32614 12939 32666
rect 12939 32614 12953 32666
rect 12977 32614 12991 32666
rect 12991 32614 13003 32666
rect 13003 32614 13033 32666
rect 13057 32614 13067 32666
rect 13067 32614 13113 32666
rect 12817 32612 12873 32614
rect 12897 32612 12953 32614
rect 12977 32612 13033 32614
rect 13057 32612 13113 32614
rect 12817 31578 12873 31580
rect 12897 31578 12953 31580
rect 12977 31578 13033 31580
rect 13057 31578 13113 31580
rect 12817 31526 12863 31578
rect 12863 31526 12873 31578
rect 12897 31526 12927 31578
rect 12927 31526 12939 31578
rect 12939 31526 12953 31578
rect 12977 31526 12991 31578
rect 12991 31526 13003 31578
rect 13003 31526 13033 31578
rect 13057 31526 13067 31578
rect 13067 31526 13113 31578
rect 12817 31524 12873 31526
rect 12897 31524 12953 31526
rect 12977 31524 13033 31526
rect 13057 31524 13113 31526
rect 3921 31034 3977 31036
rect 4001 31034 4057 31036
rect 4081 31034 4137 31036
rect 4161 31034 4217 31036
rect 3921 30982 3967 31034
rect 3967 30982 3977 31034
rect 4001 30982 4031 31034
rect 4031 30982 4043 31034
rect 4043 30982 4057 31034
rect 4081 30982 4095 31034
rect 4095 30982 4107 31034
rect 4107 30982 4137 31034
rect 4161 30982 4171 31034
rect 4171 30982 4217 31034
rect 3921 30980 3977 30982
rect 4001 30980 4057 30982
rect 4081 30980 4137 30982
rect 4161 30980 4217 30982
rect 9852 31034 9908 31036
rect 9932 31034 9988 31036
rect 10012 31034 10068 31036
rect 10092 31034 10148 31036
rect 9852 30982 9898 31034
rect 9898 30982 9908 31034
rect 9932 30982 9962 31034
rect 9962 30982 9974 31034
rect 9974 30982 9988 31034
rect 10012 30982 10026 31034
rect 10026 30982 10038 31034
rect 10038 30982 10068 31034
rect 10092 30982 10102 31034
rect 10102 30982 10148 31034
rect 9852 30980 9908 30982
rect 9932 30980 9988 30982
rect 10012 30980 10068 30982
rect 10092 30980 10148 30982
rect 1398 30504 1454 30560
rect 6886 30490 6942 30492
rect 6966 30490 7022 30492
rect 7046 30490 7102 30492
rect 7126 30490 7182 30492
rect 6886 30438 6932 30490
rect 6932 30438 6942 30490
rect 6966 30438 6996 30490
rect 6996 30438 7008 30490
rect 7008 30438 7022 30490
rect 7046 30438 7060 30490
rect 7060 30438 7072 30490
rect 7072 30438 7102 30490
rect 7126 30438 7136 30490
rect 7136 30438 7182 30490
rect 6886 30436 6942 30438
rect 6966 30436 7022 30438
rect 7046 30436 7102 30438
rect 7126 30436 7182 30438
rect 3921 29946 3977 29948
rect 4001 29946 4057 29948
rect 4081 29946 4137 29948
rect 4161 29946 4217 29948
rect 3921 29894 3967 29946
rect 3967 29894 3977 29946
rect 4001 29894 4031 29946
rect 4031 29894 4043 29946
rect 4043 29894 4057 29946
rect 4081 29894 4095 29946
rect 4095 29894 4107 29946
rect 4107 29894 4137 29946
rect 4161 29894 4171 29946
rect 4171 29894 4217 29946
rect 3921 29892 3977 29894
rect 4001 29892 4057 29894
rect 4081 29892 4137 29894
rect 4161 29892 4217 29894
rect 9852 29946 9908 29948
rect 9932 29946 9988 29948
rect 10012 29946 10068 29948
rect 10092 29946 10148 29948
rect 9852 29894 9898 29946
rect 9898 29894 9908 29946
rect 9932 29894 9962 29946
rect 9962 29894 9974 29946
rect 9974 29894 9988 29946
rect 10012 29894 10026 29946
rect 10026 29894 10038 29946
rect 10038 29894 10068 29946
rect 10092 29894 10102 29946
rect 10102 29894 10148 29946
rect 9852 29892 9908 29894
rect 9932 29892 9988 29894
rect 10012 29892 10068 29894
rect 10092 29892 10148 29894
rect 6886 29402 6942 29404
rect 6966 29402 7022 29404
rect 7046 29402 7102 29404
rect 7126 29402 7182 29404
rect 6886 29350 6932 29402
rect 6932 29350 6942 29402
rect 6966 29350 6996 29402
rect 6996 29350 7008 29402
rect 7008 29350 7022 29402
rect 7046 29350 7060 29402
rect 7060 29350 7072 29402
rect 7072 29350 7102 29402
rect 7126 29350 7136 29402
rect 7136 29350 7182 29402
rect 6886 29348 6942 29350
rect 6966 29348 7022 29350
rect 7046 29348 7102 29350
rect 7126 29348 7182 29350
rect 3921 28858 3977 28860
rect 4001 28858 4057 28860
rect 4081 28858 4137 28860
rect 4161 28858 4217 28860
rect 3921 28806 3967 28858
rect 3967 28806 3977 28858
rect 4001 28806 4031 28858
rect 4031 28806 4043 28858
rect 4043 28806 4057 28858
rect 4081 28806 4095 28858
rect 4095 28806 4107 28858
rect 4107 28806 4137 28858
rect 4161 28806 4171 28858
rect 4171 28806 4217 28858
rect 3921 28804 3977 28806
rect 4001 28804 4057 28806
rect 4081 28804 4137 28806
rect 4161 28804 4217 28806
rect 9852 28858 9908 28860
rect 9932 28858 9988 28860
rect 10012 28858 10068 28860
rect 10092 28858 10148 28860
rect 9852 28806 9898 28858
rect 9898 28806 9908 28858
rect 9932 28806 9962 28858
rect 9962 28806 9974 28858
rect 9974 28806 9988 28858
rect 10012 28806 10026 28858
rect 10026 28806 10038 28858
rect 10038 28806 10068 28858
rect 10092 28806 10102 28858
rect 10102 28806 10148 28858
rect 9852 28804 9908 28806
rect 9932 28804 9988 28806
rect 10012 28804 10068 28806
rect 10092 28804 10148 28806
rect 6886 28314 6942 28316
rect 6966 28314 7022 28316
rect 7046 28314 7102 28316
rect 7126 28314 7182 28316
rect 6886 28262 6932 28314
rect 6932 28262 6942 28314
rect 6966 28262 6996 28314
rect 6996 28262 7008 28314
rect 7008 28262 7022 28314
rect 7046 28262 7060 28314
rect 7060 28262 7072 28314
rect 7072 28262 7102 28314
rect 7126 28262 7136 28314
rect 7136 28262 7182 28314
rect 6886 28260 6942 28262
rect 6966 28260 7022 28262
rect 7046 28260 7102 28262
rect 7126 28260 7182 28262
rect 3921 27770 3977 27772
rect 4001 27770 4057 27772
rect 4081 27770 4137 27772
rect 4161 27770 4217 27772
rect 3921 27718 3967 27770
rect 3967 27718 3977 27770
rect 4001 27718 4031 27770
rect 4031 27718 4043 27770
rect 4043 27718 4057 27770
rect 4081 27718 4095 27770
rect 4095 27718 4107 27770
rect 4107 27718 4137 27770
rect 4161 27718 4171 27770
rect 4171 27718 4217 27770
rect 3921 27716 3977 27718
rect 4001 27716 4057 27718
rect 4081 27716 4137 27718
rect 4161 27716 4217 27718
rect 9852 27770 9908 27772
rect 9932 27770 9988 27772
rect 10012 27770 10068 27772
rect 10092 27770 10148 27772
rect 9852 27718 9898 27770
rect 9898 27718 9908 27770
rect 9932 27718 9962 27770
rect 9962 27718 9974 27770
rect 9974 27718 9988 27770
rect 10012 27718 10026 27770
rect 10026 27718 10038 27770
rect 10038 27718 10068 27770
rect 10092 27718 10102 27770
rect 10102 27718 10148 27770
rect 9852 27716 9908 27718
rect 9932 27716 9988 27718
rect 10012 27716 10068 27718
rect 10092 27716 10148 27718
rect 6886 27226 6942 27228
rect 6966 27226 7022 27228
rect 7046 27226 7102 27228
rect 7126 27226 7182 27228
rect 6886 27174 6932 27226
rect 6932 27174 6942 27226
rect 6966 27174 6996 27226
rect 6996 27174 7008 27226
rect 7008 27174 7022 27226
rect 7046 27174 7060 27226
rect 7060 27174 7072 27226
rect 7072 27174 7102 27226
rect 7126 27174 7136 27226
rect 7136 27174 7182 27226
rect 6886 27172 6942 27174
rect 6966 27172 7022 27174
rect 7046 27172 7102 27174
rect 7126 27172 7182 27174
rect 3921 26682 3977 26684
rect 4001 26682 4057 26684
rect 4081 26682 4137 26684
rect 4161 26682 4217 26684
rect 3921 26630 3967 26682
rect 3967 26630 3977 26682
rect 4001 26630 4031 26682
rect 4031 26630 4043 26682
rect 4043 26630 4057 26682
rect 4081 26630 4095 26682
rect 4095 26630 4107 26682
rect 4107 26630 4137 26682
rect 4161 26630 4171 26682
rect 4171 26630 4217 26682
rect 3921 26628 3977 26630
rect 4001 26628 4057 26630
rect 4081 26628 4137 26630
rect 4161 26628 4217 26630
rect 9852 26682 9908 26684
rect 9932 26682 9988 26684
rect 10012 26682 10068 26684
rect 10092 26682 10148 26684
rect 9852 26630 9898 26682
rect 9898 26630 9908 26682
rect 9932 26630 9962 26682
rect 9962 26630 9974 26682
rect 9974 26630 9988 26682
rect 10012 26630 10026 26682
rect 10026 26630 10038 26682
rect 10038 26630 10068 26682
rect 10092 26630 10102 26682
rect 10102 26630 10148 26682
rect 9852 26628 9908 26630
rect 9932 26628 9988 26630
rect 10012 26628 10068 26630
rect 10092 26628 10148 26630
rect 6886 26138 6942 26140
rect 6966 26138 7022 26140
rect 7046 26138 7102 26140
rect 7126 26138 7182 26140
rect 6886 26086 6932 26138
rect 6932 26086 6942 26138
rect 6966 26086 6996 26138
rect 6996 26086 7008 26138
rect 7008 26086 7022 26138
rect 7046 26086 7060 26138
rect 7060 26086 7072 26138
rect 7072 26086 7102 26138
rect 7126 26086 7136 26138
rect 7136 26086 7182 26138
rect 6886 26084 6942 26086
rect 6966 26084 7022 26086
rect 7046 26084 7102 26086
rect 7126 26084 7182 26086
rect 3921 25594 3977 25596
rect 4001 25594 4057 25596
rect 4081 25594 4137 25596
rect 4161 25594 4217 25596
rect 3921 25542 3967 25594
rect 3967 25542 3977 25594
rect 4001 25542 4031 25594
rect 4031 25542 4043 25594
rect 4043 25542 4057 25594
rect 4081 25542 4095 25594
rect 4095 25542 4107 25594
rect 4107 25542 4137 25594
rect 4161 25542 4171 25594
rect 4171 25542 4217 25594
rect 3921 25540 3977 25542
rect 4001 25540 4057 25542
rect 4081 25540 4137 25542
rect 4161 25540 4217 25542
rect 9852 25594 9908 25596
rect 9932 25594 9988 25596
rect 10012 25594 10068 25596
rect 10092 25594 10148 25596
rect 9852 25542 9898 25594
rect 9898 25542 9908 25594
rect 9932 25542 9962 25594
rect 9962 25542 9974 25594
rect 9974 25542 9988 25594
rect 10012 25542 10026 25594
rect 10026 25542 10038 25594
rect 10038 25542 10068 25594
rect 10092 25542 10102 25594
rect 10102 25542 10148 25594
rect 9852 25540 9908 25542
rect 9932 25540 9988 25542
rect 10012 25540 10068 25542
rect 10092 25540 10148 25542
rect 6886 25050 6942 25052
rect 6966 25050 7022 25052
rect 7046 25050 7102 25052
rect 7126 25050 7182 25052
rect 6886 24998 6932 25050
rect 6932 24998 6942 25050
rect 6966 24998 6996 25050
rect 6996 24998 7008 25050
rect 7008 24998 7022 25050
rect 7046 24998 7060 25050
rect 7060 24998 7072 25050
rect 7072 24998 7102 25050
rect 7126 24998 7136 25050
rect 7136 24998 7182 25050
rect 6886 24996 6942 24998
rect 6966 24996 7022 24998
rect 7046 24996 7102 24998
rect 7126 24996 7182 24998
rect 1490 24928 1546 24984
rect 3921 24506 3977 24508
rect 4001 24506 4057 24508
rect 4081 24506 4137 24508
rect 4161 24506 4217 24508
rect 3921 24454 3967 24506
rect 3967 24454 3977 24506
rect 4001 24454 4031 24506
rect 4031 24454 4043 24506
rect 4043 24454 4057 24506
rect 4081 24454 4095 24506
rect 4095 24454 4107 24506
rect 4107 24454 4137 24506
rect 4161 24454 4171 24506
rect 4171 24454 4217 24506
rect 3921 24452 3977 24454
rect 4001 24452 4057 24454
rect 4081 24452 4137 24454
rect 4161 24452 4217 24454
rect 9852 24506 9908 24508
rect 9932 24506 9988 24508
rect 10012 24506 10068 24508
rect 10092 24506 10148 24508
rect 9852 24454 9898 24506
rect 9898 24454 9908 24506
rect 9932 24454 9962 24506
rect 9962 24454 9974 24506
rect 9974 24454 9988 24506
rect 10012 24454 10026 24506
rect 10026 24454 10038 24506
rect 10038 24454 10068 24506
rect 10092 24454 10102 24506
rect 10102 24454 10148 24506
rect 9852 24452 9908 24454
rect 9932 24452 9988 24454
rect 10012 24452 10068 24454
rect 10092 24452 10148 24454
rect 6886 23962 6942 23964
rect 6966 23962 7022 23964
rect 7046 23962 7102 23964
rect 7126 23962 7182 23964
rect 6886 23910 6932 23962
rect 6932 23910 6942 23962
rect 6966 23910 6996 23962
rect 6996 23910 7008 23962
rect 7008 23910 7022 23962
rect 7046 23910 7060 23962
rect 7060 23910 7072 23962
rect 7072 23910 7102 23962
rect 7126 23910 7136 23962
rect 7136 23910 7182 23962
rect 6886 23908 6942 23910
rect 6966 23908 7022 23910
rect 7046 23908 7102 23910
rect 7126 23908 7182 23910
rect 3921 23418 3977 23420
rect 4001 23418 4057 23420
rect 4081 23418 4137 23420
rect 4161 23418 4217 23420
rect 3921 23366 3967 23418
rect 3967 23366 3977 23418
rect 4001 23366 4031 23418
rect 4031 23366 4043 23418
rect 4043 23366 4057 23418
rect 4081 23366 4095 23418
rect 4095 23366 4107 23418
rect 4107 23366 4137 23418
rect 4161 23366 4171 23418
rect 4171 23366 4217 23418
rect 3921 23364 3977 23366
rect 4001 23364 4057 23366
rect 4081 23364 4137 23366
rect 4161 23364 4217 23366
rect 9852 23418 9908 23420
rect 9932 23418 9988 23420
rect 10012 23418 10068 23420
rect 10092 23418 10148 23420
rect 9852 23366 9898 23418
rect 9898 23366 9908 23418
rect 9932 23366 9962 23418
rect 9962 23366 9974 23418
rect 9974 23366 9988 23418
rect 10012 23366 10026 23418
rect 10026 23366 10038 23418
rect 10038 23366 10068 23418
rect 10092 23366 10102 23418
rect 10102 23366 10148 23418
rect 9852 23364 9908 23366
rect 9932 23364 9988 23366
rect 10012 23364 10068 23366
rect 10092 23364 10148 23366
rect 6886 22874 6942 22876
rect 6966 22874 7022 22876
rect 7046 22874 7102 22876
rect 7126 22874 7182 22876
rect 6886 22822 6932 22874
rect 6932 22822 6942 22874
rect 6966 22822 6996 22874
rect 6996 22822 7008 22874
rect 7008 22822 7022 22874
rect 7046 22822 7060 22874
rect 7060 22822 7072 22874
rect 7072 22822 7102 22874
rect 7126 22822 7136 22874
rect 7136 22822 7182 22874
rect 6886 22820 6942 22822
rect 6966 22820 7022 22822
rect 7046 22820 7102 22822
rect 7126 22820 7182 22822
rect 3921 22330 3977 22332
rect 4001 22330 4057 22332
rect 4081 22330 4137 22332
rect 4161 22330 4217 22332
rect 3921 22278 3967 22330
rect 3967 22278 3977 22330
rect 4001 22278 4031 22330
rect 4031 22278 4043 22330
rect 4043 22278 4057 22330
rect 4081 22278 4095 22330
rect 4095 22278 4107 22330
rect 4107 22278 4137 22330
rect 4161 22278 4171 22330
rect 4171 22278 4217 22330
rect 3921 22276 3977 22278
rect 4001 22276 4057 22278
rect 4081 22276 4137 22278
rect 4161 22276 4217 22278
rect 9852 22330 9908 22332
rect 9932 22330 9988 22332
rect 10012 22330 10068 22332
rect 10092 22330 10148 22332
rect 9852 22278 9898 22330
rect 9898 22278 9908 22330
rect 9932 22278 9962 22330
rect 9962 22278 9974 22330
rect 9974 22278 9988 22330
rect 10012 22278 10026 22330
rect 10026 22278 10038 22330
rect 10038 22278 10068 22330
rect 10092 22278 10102 22330
rect 10102 22278 10148 22330
rect 9852 22276 9908 22278
rect 9932 22276 9988 22278
rect 10012 22276 10068 22278
rect 10092 22276 10148 22278
rect 6886 21786 6942 21788
rect 6966 21786 7022 21788
rect 7046 21786 7102 21788
rect 7126 21786 7182 21788
rect 6886 21734 6932 21786
rect 6932 21734 6942 21786
rect 6966 21734 6996 21786
rect 6996 21734 7008 21786
rect 7008 21734 7022 21786
rect 7046 21734 7060 21786
rect 7060 21734 7072 21786
rect 7072 21734 7102 21786
rect 7126 21734 7136 21786
rect 7136 21734 7182 21786
rect 6886 21732 6942 21734
rect 6966 21732 7022 21734
rect 7046 21732 7102 21734
rect 7126 21732 7182 21734
rect 3921 21242 3977 21244
rect 4001 21242 4057 21244
rect 4081 21242 4137 21244
rect 4161 21242 4217 21244
rect 3921 21190 3967 21242
rect 3967 21190 3977 21242
rect 4001 21190 4031 21242
rect 4031 21190 4043 21242
rect 4043 21190 4057 21242
rect 4081 21190 4095 21242
rect 4095 21190 4107 21242
rect 4107 21190 4137 21242
rect 4161 21190 4171 21242
rect 4171 21190 4217 21242
rect 3921 21188 3977 21190
rect 4001 21188 4057 21190
rect 4081 21188 4137 21190
rect 4161 21188 4217 21190
rect 9852 21242 9908 21244
rect 9932 21242 9988 21244
rect 10012 21242 10068 21244
rect 10092 21242 10148 21244
rect 9852 21190 9898 21242
rect 9898 21190 9908 21242
rect 9932 21190 9962 21242
rect 9962 21190 9974 21242
rect 9974 21190 9988 21242
rect 10012 21190 10026 21242
rect 10026 21190 10038 21242
rect 10038 21190 10068 21242
rect 10092 21190 10102 21242
rect 10102 21190 10148 21242
rect 9852 21188 9908 21190
rect 9932 21188 9988 21190
rect 10012 21188 10068 21190
rect 10092 21188 10148 21190
rect 6886 20698 6942 20700
rect 6966 20698 7022 20700
rect 7046 20698 7102 20700
rect 7126 20698 7182 20700
rect 6886 20646 6932 20698
rect 6932 20646 6942 20698
rect 6966 20646 6996 20698
rect 6996 20646 7008 20698
rect 7008 20646 7022 20698
rect 7046 20646 7060 20698
rect 7060 20646 7072 20698
rect 7072 20646 7102 20698
rect 7126 20646 7136 20698
rect 7136 20646 7182 20698
rect 6886 20644 6942 20646
rect 6966 20644 7022 20646
rect 7046 20644 7102 20646
rect 7126 20644 7182 20646
rect 3921 20154 3977 20156
rect 4001 20154 4057 20156
rect 4081 20154 4137 20156
rect 4161 20154 4217 20156
rect 3921 20102 3967 20154
rect 3967 20102 3977 20154
rect 4001 20102 4031 20154
rect 4031 20102 4043 20154
rect 4043 20102 4057 20154
rect 4081 20102 4095 20154
rect 4095 20102 4107 20154
rect 4107 20102 4137 20154
rect 4161 20102 4171 20154
rect 4171 20102 4217 20154
rect 3921 20100 3977 20102
rect 4001 20100 4057 20102
rect 4081 20100 4137 20102
rect 4161 20100 4217 20102
rect 9852 20154 9908 20156
rect 9932 20154 9988 20156
rect 10012 20154 10068 20156
rect 10092 20154 10148 20156
rect 9852 20102 9898 20154
rect 9898 20102 9908 20154
rect 9932 20102 9962 20154
rect 9962 20102 9974 20154
rect 9974 20102 9988 20154
rect 10012 20102 10026 20154
rect 10026 20102 10038 20154
rect 10038 20102 10068 20154
rect 10092 20102 10102 20154
rect 10102 20102 10148 20154
rect 9852 20100 9908 20102
rect 9932 20100 9988 20102
rect 10012 20100 10068 20102
rect 10092 20100 10148 20102
rect 6886 19610 6942 19612
rect 6966 19610 7022 19612
rect 7046 19610 7102 19612
rect 7126 19610 7182 19612
rect 6886 19558 6932 19610
rect 6932 19558 6942 19610
rect 6966 19558 6996 19610
rect 6996 19558 7008 19610
rect 7008 19558 7022 19610
rect 7046 19558 7060 19610
rect 7060 19558 7072 19610
rect 7072 19558 7102 19610
rect 7126 19558 7136 19610
rect 7136 19558 7182 19610
rect 6886 19556 6942 19558
rect 6966 19556 7022 19558
rect 7046 19556 7102 19558
rect 7126 19556 7182 19558
rect 1398 19388 1400 19408
rect 1400 19388 1452 19408
rect 1452 19388 1454 19408
rect 1398 19352 1454 19388
rect 3921 19066 3977 19068
rect 4001 19066 4057 19068
rect 4081 19066 4137 19068
rect 4161 19066 4217 19068
rect 3921 19014 3967 19066
rect 3967 19014 3977 19066
rect 4001 19014 4031 19066
rect 4031 19014 4043 19066
rect 4043 19014 4057 19066
rect 4081 19014 4095 19066
rect 4095 19014 4107 19066
rect 4107 19014 4137 19066
rect 4161 19014 4171 19066
rect 4171 19014 4217 19066
rect 3921 19012 3977 19014
rect 4001 19012 4057 19014
rect 4081 19012 4137 19014
rect 4161 19012 4217 19014
rect 9852 19066 9908 19068
rect 9932 19066 9988 19068
rect 10012 19066 10068 19068
rect 10092 19066 10148 19068
rect 9852 19014 9898 19066
rect 9898 19014 9908 19066
rect 9932 19014 9962 19066
rect 9962 19014 9974 19066
rect 9974 19014 9988 19066
rect 10012 19014 10026 19066
rect 10026 19014 10038 19066
rect 10038 19014 10068 19066
rect 10092 19014 10102 19066
rect 10102 19014 10148 19066
rect 9852 19012 9908 19014
rect 9932 19012 9988 19014
rect 10012 19012 10068 19014
rect 10092 19012 10148 19014
rect 6886 18522 6942 18524
rect 6966 18522 7022 18524
rect 7046 18522 7102 18524
rect 7126 18522 7182 18524
rect 6886 18470 6932 18522
rect 6932 18470 6942 18522
rect 6966 18470 6996 18522
rect 6996 18470 7008 18522
rect 7008 18470 7022 18522
rect 7046 18470 7060 18522
rect 7060 18470 7072 18522
rect 7072 18470 7102 18522
rect 7126 18470 7136 18522
rect 7136 18470 7182 18522
rect 6886 18468 6942 18470
rect 6966 18468 7022 18470
rect 7046 18468 7102 18470
rect 7126 18468 7182 18470
rect 3921 17978 3977 17980
rect 4001 17978 4057 17980
rect 4081 17978 4137 17980
rect 4161 17978 4217 17980
rect 3921 17926 3967 17978
rect 3967 17926 3977 17978
rect 4001 17926 4031 17978
rect 4031 17926 4043 17978
rect 4043 17926 4057 17978
rect 4081 17926 4095 17978
rect 4095 17926 4107 17978
rect 4107 17926 4137 17978
rect 4161 17926 4171 17978
rect 4171 17926 4217 17978
rect 3921 17924 3977 17926
rect 4001 17924 4057 17926
rect 4081 17924 4137 17926
rect 4161 17924 4217 17926
rect 6886 17434 6942 17436
rect 6966 17434 7022 17436
rect 7046 17434 7102 17436
rect 7126 17434 7182 17436
rect 6886 17382 6932 17434
rect 6932 17382 6942 17434
rect 6966 17382 6996 17434
rect 6996 17382 7008 17434
rect 7008 17382 7022 17434
rect 7046 17382 7060 17434
rect 7060 17382 7072 17434
rect 7072 17382 7102 17434
rect 7126 17382 7136 17434
rect 7136 17382 7182 17434
rect 6886 17380 6942 17382
rect 6966 17380 7022 17382
rect 7046 17380 7102 17382
rect 7126 17380 7182 17382
rect 3921 16890 3977 16892
rect 4001 16890 4057 16892
rect 4081 16890 4137 16892
rect 4161 16890 4217 16892
rect 3921 16838 3967 16890
rect 3967 16838 3977 16890
rect 4001 16838 4031 16890
rect 4031 16838 4043 16890
rect 4043 16838 4057 16890
rect 4081 16838 4095 16890
rect 4095 16838 4107 16890
rect 4107 16838 4137 16890
rect 4161 16838 4171 16890
rect 4171 16838 4217 16890
rect 3921 16836 3977 16838
rect 4001 16836 4057 16838
rect 4081 16836 4137 16838
rect 4161 16836 4217 16838
rect 6886 16346 6942 16348
rect 6966 16346 7022 16348
rect 7046 16346 7102 16348
rect 7126 16346 7182 16348
rect 6886 16294 6932 16346
rect 6932 16294 6942 16346
rect 6966 16294 6996 16346
rect 6996 16294 7008 16346
rect 7008 16294 7022 16346
rect 7046 16294 7060 16346
rect 7060 16294 7072 16346
rect 7072 16294 7102 16346
rect 7126 16294 7136 16346
rect 7136 16294 7182 16346
rect 6886 16292 6942 16294
rect 6966 16292 7022 16294
rect 7046 16292 7102 16294
rect 7126 16292 7182 16294
rect 3921 15802 3977 15804
rect 4001 15802 4057 15804
rect 4081 15802 4137 15804
rect 4161 15802 4217 15804
rect 3921 15750 3967 15802
rect 3967 15750 3977 15802
rect 4001 15750 4031 15802
rect 4031 15750 4043 15802
rect 4043 15750 4057 15802
rect 4081 15750 4095 15802
rect 4095 15750 4107 15802
rect 4107 15750 4137 15802
rect 4161 15750 4171 15802
rect 4171 15750 4217 15802
rect 3921 15748 3977 15750
rect 4001 15748 4057 15750
rect 4081 15748 4137 15750
rect 4161 15748 4217 15750
rect 6886 15258 6942 15260
rect 6966 15258 7022 15260
rect 7046 15258 7102 15260
rect 7126 15258 7182 15260
rect 6886 15206 6932 15258
rect 6932 15206 6942 15258
rect 6966 15206 6996 15258
rect 6996 15206 7008 15258
rect 7008 15206 7022 15258
rect 7046 15206 7060 15258
rect 7060 15206 7072 15258
rect 7072 15206 7102 15258
rect 7126 15206 7136 15258
rect 7136 15206 7182 15258
rect 6886 15204 6942 15206
rect 6966 15204 7022 15206
rect 7046 15204 7102 15206
rect 7126 15204 7182 15206
rect 3921 14714 3977 14716
rect 4001 14714 4057 14716
rect 4081 14714 4137 14716
rect 4161 14714 4217 14716
rect 3921 14662 3967 14714
rect 3967 14662 3977 14714
rect 4001 14662 4031 14714
rect 4031 14662 4043 14714
rect 4043 14662 4057 14714
rect 4081 14662 4095 14714
rect 4095 14662 4107 14714
rect 4107 14662 4137 14714
rect 4161 14662 4171 14714
rect 4171 14662 4217 14714
rect 3921 14660 3977 14662
rect 4001 14660 4057 14662
rect 4081 14660 4137 14662
rect 4161 14660 4217 14662
rect 6886 14170 6942 14172
rect 6966 14170 7022 14172
rect 7046 14170 7102 14172
rect 7126 14170 7182 14172
rect 6886 14118 6932 14170
rect 6932 14118 6942 14170
rect 6966 14118 6996 14170
rect 6996 14118 7008 14170
rect 7008 14118 7022 14170
rect 7046 14118 7060 14170
rect 7060 14118 7072 14170
rect 7072 14118 7102 14170
rect 7126 14118 7136 14170
rect 7136 14118 7182 14170
rect 6886 14116 6942 14118
rect 6966 14116 7022 14118
rect 7046 14116 7102 14118
rect 7126 14116 7182 14118
rect 9852 17978 9908 17980
rect 9932 17978 9988 17980
rect 10012 17978 10068 17980
rect 10092 17978 10148 17980
rect 9852 17926 9898 17978
rect 9898 17926 9908 17978
rect 9932 17926 9962 17978
rect 9962 17926 9974 17978
rect 9974 17926 9988 17978
rect 10012 17926 10026 17978
rect 10026 17926 10038 17978
rect 10038 17926 10068 17978
rect 10092 17926 10102 17978
rect 10102 17926 10148 17978
rect 9852 17924 9908 17926
rect 9932 17924 9988 17926
rect 10012 17924 10068 17926
rect 10092 17924 10148 17926
rect 9852 16890 9908 16892
rect 9932 16890 9988 16892
rect 10012 16890 10068 16892
rect 10092 16890 10148 16892
rect 9852 16838 9898 16890
rect 9898 16838 9908 16890
rect 9932 16838 9962 16890
rect 9962 16838 9974 16890
rect 9974 16838 9988 16890
rect 10012 16838 10026 16890
rect 10026 16838 10038 16890
rect 10038 16838 10068 16890
rect 10092 16838 10102 16890
rect 10102 16838 10148 16890
rect 9852 16836 9908 16838
rect 9932 16836 9988 16838
rect 10012 16836 10068 16838
rect 10092 16836 10148 16838
rect 9852 15802 9908 15804
rect 9932 15802 9988 15804
rect 10012 15802 10068 15804
rect 10092 15802 10148 15804
rect 9852 15750 9898 15802
rect 9898 15750 9908 15802
rect 9932 15750 9962 15802
rect 9962 15750 9974 15802
rect 9974 15750 9988 15802
rect 10012 15750 10026 15802
rect 10026 15750 10038 15802
rect 10038 15750 10068 15802
rect 10092 15750 10102 15802
rect 10102 15750 10148 15802
rect 9852 15748 9908 15750
rect 9932 15748 9988 15750
rect 10012 15748 10068 15750
rect 10092 15748 10148 15750
rect 9852 14714 9908 14716
rect 9932 14714 9988 14716
rect 10012 14714 10068 14716
rect 10092 14714 10148 14716
rect 9852 14662 9898 14714
rect 9898 14662 9908 14714
rect 9932 14662 9962 14714
rect 9962 14662 9974 14714
rect 9974 14662 9988 14714
rect 10012 14662 10026 14714
rect 10026 14662 10038 14714
rect 10038 14662 10068 14714
rect 10092 14662 10102 14714
rect 10102 14662 10148 14714
rect 9852 14660 9908 14662
rect 9932 14660 9988 14662
rect 10012 14660 10068 14662
rect 10092 14660 10148 14662
rect 1398 13812 1400 13832
rect 1400 13812 1452 13832
rect 1452 13812 1454 13832
rect 1398 13776 1454 13812
rect 3921 13626 3977 13628
rect 4001 13626 4057 13628
rect 4081 13626 4137 13628
rect 4161 13626 4217 13628
rect 3921 13574 3967 13626
rect 3967 13574 3977 13626
rect 4001 13574 4031 13626
rect 4031 13574 4043 13626
rect 4043 13574 4057 13626
rect 4081 13574 4095 13626
rect 4095 13574 4107 13626
rect 4107 13574 4137 13626
rect 4161 13574 4171 13626
rect 4171 13574 4217 13626
rect 3921 13572 3977 13574
rect 4001 13572 4057 13574
rect 4081 13572 4137 13574
rect 4161 13572 4217 13574
rect 9852 13626 9908 13628
rect 9932 13626 9988 13628
rect 10012 13626 10068 13628
rect 10092 13626 10148 13628
rect 9852 13574 9898 13626
rect 9898 13574 9908 13626
rect 9932 13574 9962 13626
rect 9962 13574 9974 13626
rect 9974 13574 9988 13626
rect 10012 13574 10026 13626
rect 10026 13574 10038 13626
rect 10038 13574 10068 13626
rect 10092 13574 10102 13626
rect 10102 13574 10148 13626
rect 9852 13572 9908 13574
rect 9932 13572 9988 13574
rect 10012 13572 10068 13574
rect 10092 13572 10148 13574
rect 6886 13082 6942 13084
rect 6966 13082 7022 13084
rect 7046 13082 7102 13084
rect 7126 13082 7182 13084
rect 6886 13030 6932 13082
rect 6932 13030 6942 13082
rect 6966 13030 6996 13082
rect 6996 13030 7008 13082
rect 7008 13030 7022 13082
rect 7046 13030 7060 13082
rect 7060 13030 7072 13082
rect 7072 13030 7102 13082
rect 7126 13030 7136 13082
rect 7136 13030 7182 13082
rect 6886 13028 6942 13030
rect 6966 13028 7022 13030
rect 7046 13028 7102 13030
rect 7126 13028 7182 13030
rect 3921 12538 3977 12540
rect 4001 12538 4057 12540
rect 4081 12538 4137 12540
rect 4161 12538 4217 12540
rect 3921 12486 3967 12538
rect 3967 12486 3977 12538
rect 4001 12486 4031 12538
rect 4031 12486 4043 12538
rect 4043 12486 4057 12538
rect 4081 12486 4095 12538
rect 4095 12486 4107 12538
rect 4107 12486 4137 12538
rect 4161 12486 4171 12538
rect 4171 12486 4217 12538
rect 3921 12484 3977 12486
rect 4001 12484 4057 12486
rect 4081 12484 4137 12486
rect 4161 12484 4217 12486
rect 9852 12538 9908 12540
rect 9932 12538 9988 12540
rect 10012 12538 10068 12540
rect 10092 12538 10148 12540
rect 9852 12486 9898 12538
rect 9898 12486 9908 12538
rect 9932 12486 9962 12538
rect 9962 12486 9974 12538
rect 9974 12486 9988 12538
rect 10012 12486 10026 12538
rect 10026 12486 10038 12538
rect 10038 12486 10068 12538
rect 10092 12486 10102 12538
rect 10102 12486 10148 12538
rect 9852 12484 9908 12486
rect 9932 12484 9988 12486
rect 10012 12484 10068 12486
rect 10092 12484 10148 12486
rect 6886 11994 6942 11996
rect 6966 11994 7022 11996
rect 7046 11994 7102 11996
rect 7126 11994 7182 11996
rect 6886 11942 6932 11994
rect 6932 11942 6942 11994
rect 6966 11942 6996 11994
rect 6996 11942 7008 11994
rect 7008 11942 7022 11994
rect 7046 11942 7060 11994
rect 7060 11942 7072 11994
rect 7072 11942 7102 11994
rect 7126 11942 7136 11994
rect 7136 11942 7182 11994
rect 6886 11940 6942 11942
rect 6966 11940 7022 11942
rect 7046 11940 7102 11942
rect 7126 11940 7182 11942
rect 3921 11450 3977 11452
rect 4001 11450 4057 11452
rect 4081 11450 4137 11452
rect 4161 11450 4217 11452
rect 3921 11398 3967 11450
rect 3967 11398 3977 11450
rect 4001 11398 4031 11450
rect 4031 11398 4043 11450
rect 4043 11398 4057 11450
rect 4081 11398 4095 11450
rect 4095 11398 4107 11450
rect 4107 11398 4137 11450
rect 4161 11398 4171 11450
rect 4171 11398 4217 11450
rect 3921 11396 3977 11398
rect 4001 11396 4057 11398
rect 4081 11396 4137 11398
rect 4161 11396 4217 11398
rect 9852 11450 9908 11452
rect 9932 11450 9988 11452
rect 10012 11450 10068 11452
rect 10092 11450 10148 11452
rect 9852 11398 9898 11450
rect 9898 11398 9908 11450
rect 9932 11398 9962 11450
rect 9962 11398 9974 11450
rect 9974 11398 9988 11450
rect 10012 11398 10026 11450
rect 10026 11398 10038 11450
rect 10038 11398 10068 11450
rect 10092 11398 10102 11450
rect 10102 11398 10148 11450
rect 9852 11396 9908 11398
rect 9932 11396 9988 11398
rect 10012 11396 10068 11398
rect 10092 11396 10148 11398
rect 6886 10906 6942 10908
rect 6966 10906 7022 10908
rect 7046 10906 7102 10908
rect 7126 10906 7182 10908
rect 6886 10854 6932 10906
rect 6932 10854 6942 10906
rect 6966 10854 6996 10906
rect 6996 10854 7008 10906
rect 7008 10854 7022 10906
rect 7046 10854 7060 10906
rect 7060 10854 7072 10906
rect 7072 10854 7102 10906
rect 7126 10854 7136 10906
rect 7136 10854 7182 10906
rect 6886 10852 6942 10854
rect 6966 10852 7022 10854
rect 7046 10852 7102 10854
rect 7126 10852 7182 10854
rect 3921 10362 3977 10364
rect 4001 10362 4057 10364
rect 4081 10362 4137 10364
rect 4161 10362 4217 10364
rect 3921 10310 3967 10362
rect 3967 10310 3977 10362
rect 4001 10310 4031 10362
rect 4031 10310 4043 10362
rect 4043 10310 4057 10362
rect 4081 10310 4095 10362
rect 4095 10310 4107 10362
rect 4107 10310 4137 10362
rect 4161 10310 4171 10362
rect 4171 10310 4217 10362
rect 3921 10308 3977 10310
rect 4001 10308 4057 10310
rect 4081 10308 4137 10310
rect 4161 10308 4217 10310
rect 9852 10362 9908 10364
rect 9932 10362 9988 10364
rect 10012 10362 10068 10364
rect 10092 10362 10148 10364
rect 9852 10310 9898 10362
rect 9898 10310 9908 10362
rect 9932 10310 9962 10362
rect 9962 10310 9974 10362
rect 9974 10310 9988 10362
rect 10012 10310 10026 10362
rect 10026 10310 10038 10362
rect 10038 10310 10068 10362
rect 10092 10310 10102 10362
rect 10102 10310 10148 10362
rect 9852 10308 9908 10310
rect 9932 10308 9988 10310
rect 10012 10308 10068 10310
rect 10092 10308 10148 10310
rect 6886 9818 6942 9820
rect 6966 9818 7022 9820
rect 7046 9818 7102 9820
rect 7126 9818 7182 9820
rect 6886 9766 6932 9818
rect 6932 9766 6942 9818
rect 6966 9766 6996 9818
rect 6996 9766 7008 9818
rect 7008 9766 7022 9818
rect 7046 9766 7060 9818
rect 7060 9766 7072 9818
rect 7072 9766 7102 9818
rect 7126 9766 7136 9818
rect 7136 9766 7182 9818
rect 6886 9764 6942 9766
rect 6966 9764 7022 9766
rect 7046 9764 7102 9766
rect 7126 9764 7182 9766
rect 3921 9274 3977 9276
rect 4001 9274 4057 9276
rect 4081 9274 4137 9276
rect 4161 9274 4217 9276
rect 3921 9222 3967 9274
rect 3967 9222 3977 9274
rect 4001 9222 4031 9274
rect 4031 9222 4043 9274
rect 4043 9222 4057 9274
rect 4081 9222 4095 9274
rect 4095 9222 4107 9274
rect 4107 9222 4137 9274
rect 4161 9222 4171 9274
rect 4171 9222 4217 9274
rect 3921 9220 3977 9222
rect 4001 9220 4057 9222
rect 4081 9220 4137 9222
rect 4161 9220 4217 9222
rect 9852 9274 9908 9276
rect 9932 9274 9988 9276
rect 10012 9274 10068 9276
rect 10092 9274 10148 9276
rect 9852 9222 9898 9274
rect 9898 9222 9908 9274
rect 9932 9222 9962 9274
rect 9962 9222 9974 9274
rect 9974 9222 9988 9274
rect 10012 9222 10026 9274
rect 10026 9222 10038 9274
rect 10038 9222 10068 9274
rect 10092 9222 10102 9274
rect 10102 9222 10148 9274
rect 9852 9220 9908 9222
rect 9932 9220 9988 9222
rect 10012 9220 10068 9222
rect 10092 9220 10148 9222
rect 6886 8730 6942 8732
rect 6966 8730 7022 8732
rect 7046 8730 7102 8732
rect 7126 8730 7182 8732
rect 6886 8678 6932 8730
rect 6932 8678 6942 8730
rect 6966 8678 6996 8730
rect 6996 8678 7008 8730
rect 7008 8678 7022 8730
rect 7046 8678 7060 8730
rect 7060 8678 7072 8730
rect 7072 8678 7102 8730
rect 7126 8678 7136 8730
rect 7136 8678 7182 8730
rect 6886 8676 6942 8678
rect 6966 8676 7022 8678
rect 7046 8676 7102 8678
rect 7126 8676 7182 8678
rect 1582 8200 1638 8256
rect 3921 8186 3977 8188
rect 4001 8186 4057 8188
rect 4081 8186 4137 8188
rect 4161 8186 4217 8188
rect 3921 8134 3967 8186
rect 3967 8134 3977 8186
rect 4001 8134 4031 8186
rect 4031 8134 4043 8186
rect 4043 8134 4057 8186
rect 4081 8134 4095 8186
rect 4095 8134 4107 8186
rect 4107 8134 4137 8186
rect 4161 8134 4171 8186
rect 4171 8134 4217 8186
rect 3921 8132 3977 8134
rect 4001 8132 4057 8134
rect 4081 8132 4137 8134
rect 4161 8132 4217 8134
rect 9852 8186 9908 8188
rect 9932 8186 9988 8188
rect 10012 8186 10068 8188
rect 10092 8186 10148 8188
rect 9852 8134 9898 8186
rect 9898 8134 9908 8186
rect 9932 8134 9962 8186
rect 9962 8134 9974 8186
rect 9974 8134 9988 8186
rect 10012 8134 10026 8186
rect 10026 8134 10038 8186
rect 10038 8134 10068 8186
rect 10092 8134 10102 8186
rect 10102 8134 10148 8186
rect 9852 8132 9908 8134
rect 9932 8132 9988 8134
rect 10012 8132 10068 8134
rect 10092 8132 10148 8134
rect 6886 7642 6942 7644
rect 6966 7642 7022 7644
rect 7046 7642 7102 7644
rect 7126 7642 7182 7644
rect 6886 7590 6932 7642
rect 6932 7590 6942 7642
rect 6966 7590 6996 7642
rect 6996 7590 7008 7642
rect 7008 7590 7022 7642
rect 7046 7590 7060 7642
rect 7060 7590 7072 7642
rect 7072 7590 7102 7642
rect 7126 7590 7136 7642
rect 7136 7590 7182 7642
rect 6886 7588 6942 7590
rect 6966 7588 7022 7590
rect 7046 7588 7102 7590
rect 7126 7588 7182 7590
rect 3921 7098 3977 7100
rect 4001 7098 4057 7100
rect 4081 7098 4137 7100
rect 4161 7098 4217 7100
rect 3921 7046 3967 7098
rect 3967 7046 3977 7098
rect 4001 7046 4031 7098
rect 4031 7046 4043 7098
rect 4043 7046 4057 7098
rect 4081 7046 4095 7098
rect 4095 7046 4107 7098
rect 4107 7046 4137 7098
rect 4161 7046 4171 7098
rect 4171 7046 4217 7098
rect 3921 7044 3977 7046
rect 4001 7044 4057 7046
rect 4081 7044 4137 7046
rect 4161 7044 4217 7046
rect 9852 7098 9908 7100
rect 9932 7098 9988 7100
rect 10012 7098 10068 7100
rect 10092 7098 10148 7100
rect 9852 7046 9898 7098
rect 9898 7046 9908 7098
rect 9932 7046 9962 7098
rect 9962 7046 9974 7098
rect 9974 7046 9988 7098
rect 10012 7046 10026 7098
rect 10026 7046 10038 7098
rect 10038 7046 10068 7098
rect 10092 7046 10102 7098
rect 10102 7046 10148 7098
rect 9852 7044 9908 7046
rect 9932 7044 9988 7046
rect 10012 7044 10068 7046
rect 10092 7044 10148 7046
rect 6886 6554 6942 6556
rect 6966 6554 7022 6556
rect 7046 6554 7102 6556
rect 7126 6554 7182 6556
rect 6886 6502 6932 6554
rect 6932 6502 6942 6554
rect 6966 6502 6996 6554
rect 6996 6502 7008 6554
rect 7008 6502 7022 6554
rect 7046 6502 7060 6554
rect 7060 6502 7072 6554
rect 7072 6502 7102 6554
rect 7126 6502 7136 6554
rect 7136 6502 7182 6554
rect 6886 6500 6942 6502
rect 6966 6500 7022 6502
rect 7046 6500 7102 6502
rect 7126 6500 7182 6502
rect 3921 6010 3977 6012
rect 4001 6010 4057 6012
rect 4081 6010 4137 6012
rect 4161 6010 4217 6012
rect 3921 5958 3967 6010
rect 3967 5958 3977 6010
rect 4001 5958 4031 6010
rect 4031 5958 4043 6010
rect 4043 5958 4057 6010
rect 4081 5958 4095 6010
rect 4095 5958 4107 6010
rect 4107 5958 4137 6010
rect 4161 5958 4171 6010
rect 4171 5958 4217 6010
rect 3921 5956 3977 5958
rect 4001 5956 4057 5958
rect 4081 5956 4137 5958
rect 4161 5956 4217 5958
rect 9852 6010 9908 6012
rect 9932 6010 9988 6012
rect 10012 6010 10068 6012
rect 10092 6010 10148 6012
rect 9852 5958 9898 6010
rect 9898 5958 9908 6010
rect 9932 5958 9962 6010
rect 9962 5958 9974 6010
rect 9974 5958 9988 6010
rect 10012 5958 10026 6010
rect 10026 5958 10038 6010
rect 10038 5958 10068 6010
rect 10092 5958 10102 6010
rect 10102 5958 10148 6010
rect 9852 5956 9908 5958
rect 9932 5956 9988 5958
rect 10012 5956 10068 5958
rect 10092 5956 10148 5958
rect 6886 5466 6942 5468
rect 6966 5466 7022 5468
rect 7046 5466 7102 5468
rect 7126 5466 7182 5468
rect 6886 5414 6932 5466
rect 6932 5414 6942 5466
rect 6966 5414 6996 5466
rect 6996 5414 7008 5466
rect 7008 5414 7022 5466
rect 7046 5414 7060 5466
rect 7060 5414 7072 5466
rect 7072 5414 7102 5466
rect 7126 5414 7136 5466
rect 7136 5414 7182 5466
rect 6886 5412 6942 5414
rect 6966 5412 7022 5414
rect 7046 5412 7102 5414
rect 7126 5412 7182 5414
rect 3921 4922 3977 4924
rect 4001 4922 4057 4924
rect 4081 4922 4137 4924
rect 4161 4922 4217 4924
rect 3921 4870 3967 4922
rect 3967 4870 3977 4922
rect 4001 4870 4031 4922
rect 4031 4870 4043 4922
rect 4043 4870 4057 4922
rect 4081 4870 4095 4922
rect 4095 4870 4107 4922
rect 4107 4870 4137 4922
rect 4161 4870 4171 4922
rect 4171 4870 4217 4922
rect 3921 4868 3977 4870
rect 4001 4868 4057 4870
rect 4081 4868 4137 4870
rect 4161 4868 4217 4870
rect 9852 4922 9908 4924
rect 9932 4922 9988 4924
rect 10012 4922 10068 4924
rect 10092 4922 10148 4924
rect 9852 4870 9898 4922
rect 9898 4870 9908 4922
rect 9932 4870 9962 4922
rect 9962 4870 9974 4922
rect 9974 4870 9988 4922
rect 10012 4870 10026 4922
rect 10026 4870 10038 4922
rect 10038 4870 10068 4922
rect 10092 4870 10102 4922
rect 10102 4870 10148 4922
rect 9852 4868 9908 4870
rect 9932 4868 9988 4870
rect 10012 4868 10068 4870
rect 10092 4868 10148 4870
rect 6886 4378 6942 4380
rect 6966 4378 7022 4380
rect 7046 4378 7102 4380
rect 7126 4378 7182 4380
rect 6886 4326 6932 4378
rect 6932 4326 6942 4378
rect 6966 4326 6996 4378
rect 6996 4326 7008 4378
rect 7008 4326 7022 4378
rect 7046 4326 7060 4378
rect 7060 4326 7072 4378
rect 7072 4326 7102 4378
rect 7126 4326 7136 4378
rect 7136 4326 7182 4378
rect 6886 4324 6942 4326
rect 6966 4324 7022 4326
rect 7046 4324 7102 4326
rect 7126 4324 7182 4326
rect 3921 3834 3977 3836
rect 4001 3834 4057 3836
rect 4081 3834 4137 3836
rect 4161 3834 4217 3836
rect 3921 3782 3967 3834
rect 3967 3782 3977 3834
rect 4001 3782 4031 3834
rect 4031 3782 4043 3834
rect 4043 3782 4057 3834
rect 4081 3782 4095 3834
rect 4095 3782 4107 3834
rect 4107 3782 4137 3834
rect 4161 3782 4171 3834
rect 4171 3782 4217 3834
rect 3921 3780 3977 3782
rect 4001 3780 4057 3782
rect 4081 3780 4137 3782
rect 4161 3780 4217 3782
rect 9852 3834 9908 3836
rect 9932 3834 9988 3836
rect 10012 3834 10068 3836
rect 10092 3834 10148 3836
rect 9852 3782 9898 3834
rect 9898 3782 9908 3834
rect 9932 3782 9962 3834
rect 9962 3782 9974 3834
rect 9974 3782 9988 3834
rect 10012 3782 10026 3834
rect 10026 3782 10038 3834
rect 10038 3782 10068 3834
rect 10092 3782 10102 3834
rect 10102 3782 10148 3834
rect 9852 3780 9908 3782
rect 9932 3780 9988 3782
rect 10012 3780 10068 3782
rect 10092 3780 10148 3782
rect 6886 3290 6942 3292
rect 6966 3290 7022 3292
rect 7046 3290 7102 3292
rect 7126 3290 7182 3292
rect 6886 3238 6932 3290
rect 6932 3238 6942 3290
rect 6966 3238 6996 3290
rect 6996 3238 7008 3290
rect 7008 3238 7022 3290
rect 7046 3238 7060 3290
rect 7060 3238 7072 3290
rect 7072 3238 7102 3290
rect 7126 3238 7136 3290
rect 7136 3238 7182 3290
rect 6886 3236 6942 3238
rect 6966 3236 7022 3238
rect 7046 3236 7102 3238
rect 7126 3236 7182 3238
rect 2226 2932 2228 2952
rect 2228 2932 2280 2952
rect 2280 2932 2282 2952
rect 2226 2896 2282 2932
rect 1490 2796 1492 2816
rect 1492 2796 1544 2816
rect 1544 2796 1546 2816
rect 1490 2760 1546 2796
rect 3921 2746 3977 2748
rect 4001 2746 4057 2748
rect 4081 2746 4137 2748
rect 4161 2746 4217 2748
rect 3921 2694 3967 2746
rect 3967 2694 3977 2746
rect 4001 2694 4031 2746
rect 4031 2694 4043 2746
rect 4043 2694 4057 2746
rect 4081 2694 4095 2746
rect 4095 2694 4107 2746
rect 4107 2694 4137 2746
rect 4161 2694 4171 2746
rect 4171 2694 4217 2746
rect 3921 2692 3977 2694
rect 4001 2692 4057 2694
rect 4081 2692 4137 2694
rect 4161 2692 4217 2694
rect 9852 2746 9908 2748
rect 9932 2746 9988 2748
rect 10012 2746 10068 2748
rect 10092 2746 10148 2748
rect 9852 2694 9898 2746
rect 9898 2694 9908 2746
rect 9932 2694 9962 2746
rect 9962 2694 9974 2746
rect 9974 2694 9988 2746
rect 10012 2694 10026 2746
rect 10026 2694 10038 2746
rect 10038 2694 10068 2746
rect 10092 2694 10102 2746
rect 10102 2694 10148 2746
rect 9852 2692 9908 2694
rect 9932 2692 9988 2694
rect 10012 2692 10068 2694
rect 10092 2692 10148 2694
rect 12817 30490 12873 30492
rect 12897 30490 12953 30492
rect 12977 30490 13033 30492
rect 13057 30490 13113 30492
rect 12817 30438 12863 30490
rect 12863 30438 12873 30490
rect 12897 30438 12927 30490
rect 12927 30438 12939 30490
rect 12939 30438 12953 30490
rect 12977 30438 12991 30490
rect 12991 30438 13003 30490
rect 13003 30438 13033 30490
rect 13057 30438 13067 30490
rect 13067 30438 13113 30490
rect 12817 30436 12873 30438
rect 12897 30436 12953 30438
rect 12977 30436 13033 30438
rect 13057 30436 13113 30438
rect 12817 29402 12873 29404
rect 12897 29402 12953 29404
rect 12977 29402 13033 29404
rect 13057 29402 13113 29404
rect 12817 29350 12863 29402
rect 12863 29350 12873 29402
rect 12897 29350 12927 29402
rect 12927 29350 12939 29402
rect 12939 29350 12953 29402
rect 12977 29350 12991 29402
rect 12991 29350 13003 29402
rect 13003 29350 13033 29402
rect 13057 29350 13067 29402
rect 13067 29350 13113 29402
rect 12817 29348 12873 29350
rect 12897 29348 12953 29350
rect 12977 29348 13033 29350
rect 13057 29348 13113 29350
rect 12817 28314 12873 28316
rect 12897 28314 12953 28316
rect 12977 28314 13033 28316
rect 13057 28314 13113 28316
rect 12817 28262 12863 28314
rect 12863 28262 12873 28314
rect 12897 28262 12927 28314
rect 12927 28262 12939 28314
rect 12939 28262 12953 28314
rect 12977 28262 12991 28314
rect 12991 28262 13003 28314
rect 13003 28262 13033 28314
rect 13057 28262 13067 28314
rect 13067 28262 13113 28314
rect 12817 28260 12873 28262
rect 12897 28260 12953 28262
rect 12977 28260 13033 28262
rect 13057 28260 13113 28262
rect 12817 27226 12873 27228
rect 12897 27226 12953 27228
rect 12977 27226 13033 27228
rect 13057 27226 13113 27228
rect 12817 27174 12863 27226
rect 12863 27174 12873 27226
rect 12897 27174 12927 27226
rect 12927 27174 12939 27226
rect 12939 27174 12953 27226
rect 12977 27174 12991 27226
rect 12991 27174 13003 27226
rect 13003 27174 13033 27226
rect 13057 27174 13067 27226
rect 13067 27174 13113 27226
rect 12817 27172 12873 27174
rect 12897 27172 12953 27174
rect 12977 27172 13033 27174
rect 13057 27172 13113 27174
rect 12817 26138 12873 26140
rect 12897 26138 12953 26140
rect 12977 26138 13033 26140
rect 13057 26138 13113 26140
rect 12817 26086 12863 26138
rect 12863 26086 12873 26138
rect 12897 26086 12927 26138
rect 12927 26086 12939 26138
rect 12939 26086 12953 26138
rect 12977 26086 12991 26138
rect 12991 26086 13003 26138
rect 13003 26086 13033 26138
rect 13057 26086 13067 26138
rect 13067 26086 13113 26138
rect 12817 26084 12873 26086
rect 12897 26084 12953 26086
rect 12977 26084 13033 26086
rect 13057 26084 13113 26086
rect 13174 25492 13230 25528
rect 13174 25472 13176 25492
rect 13176 25472 13228 25492
rect 13228 25472 13230 25492
rect 12817 25050 12873 25052
rect 12897 25050 12953 25052
rect 12977 25050 13033 25052
rect 13057 25050 13113 25052
rect 12817 24998 12863 25050
rect 12863 24998 12873 25050
rect 12897 24998 12927 25050
rect 12927 24998 12939 25050
rect 12939 24998 12953 25050
rect 12977 24998 12991 25050
rect 12991 24998 13003 25050
rect 13003 24998 13033 25050
rect 13057 24998 13067 25050
rect 13067 24998 13113 25050
rect 12817 24996 12873 24998
rect 12897 24996 12953 24998
rect 12977 24996 13033 24998
rect 13057 24996 13113 24998
rect 12817 23962 12873 23964
rect 12897 23962 12953 23964
rect 12977 23962 13033 23964
rect 13057 23962 13113 23964
rect 12817 23910 12863 23962
rect 12863 23910 12873 23962
rect 12897 23910 12927 23962
rect 12927 23910 12939 23962
rect 12939 23910 12953 23962
rect 12977 23910 12991 23962
rect 12991 23910 13003 23962
rect 13003 23910 13033 23962
rect 13057 23910 13067 23962
rect 13067 23910 13113 23962
rect 12817 23908 12873 23910
rect 12897 23908 12953 23910
rect 12977 23908 13033 23910
rect 13057 23908 13113 23910
rect 12817 22874 12873 22876
rect 12897 22874 12953 22876
rect 12977 22874 13033 22876
rect 13057 22874 13113 22876
rect 12817 22822 12863 22874
rect 12863 22822 12873 22874
rect 12897 22822 12927 22874
rect 12927 22822 12939 22874
rect 12939 22822 12953 22874
rect 12977 22822 12991 22874
rect 12991 22822 13003 22874
rect 13003 22822 13033 22874
rect 13057 22822 13067 22874
rect 13067 22822 13113 22874
rect 12817 22820 12873 22822
rect 12897 22820 12953 22822
rect 12977 22820 13033 22822
rect 13057 22820 13113 22822
rect 12817 21786 12873 21788
rect 12897 21786 12953 21788
rect 12977 21786 13033 21788
rect 13057 21786 13113 21788
rect 12817 21734 12863 21786
rect 12863 21734 12873 21786
rect 12897 21734 12927 21786
rect 12927 21734 12939 21786
rect 12939 21734 12953 21786
rect 12977 21734 12991 21786
rect 12991 21734 13003 21786
rect 13003 21734 13033 21786
rect 13057 21734 13067 21786
rect 13067 21734 13113 21786
rect 12817 21732 12873 21734
rect 12897 21732 12953 21734
rect 12977 21732 13033 21734
rect 13057 21732 13113 21734
rect 12817 20698 12873 20700
rect 12897 20698 12953 20700
rect 12977 20698 13033 20700
rect 13057 20698 13113 20700
rect 12817 20646 12863 20698
rect 12863 20646 12873 20698
rect 12897 20646 12927 20698
rect 12927 20646 12939 20698
rect 12939 20646 12953 20698
rect 12977 20646 12991 20698
rect 12991 20646 13003 20698
rect 13003 20646 13033 20698
rect 13057 20646 13067 20698
rect 13067 20646 13113 20698
rect 12817 20644 12873 20646
rect 12897 20644 12953 20646
rect 12977 20644 13033 20646
rect 13057 20644 13113 20646
rect 12817 19610 12873 19612
rect 12897 19610 12953 19612
rect 12977 19610 13033 19612
rect 13057 19610 13113 19612
rect 12817 19558 12863 19610
rect 12863 19558 12873 19610
rect 12897 19558 12927 19610
rect 12927 19558 12939 19610
rect 12939 19558 12953 19610
rect 12977 19558 12991 19610
rect 12991 19558 13003 19610
rect 13003 19558 13033 19610
rect 13057 19558 13067 19610
rect 13067 19558 13113 19610
rect 12817 19556 12873 19558
rect 12897 19556 12953 19558
rect 12977 19556 13033 19558
rect 13057 19556 13113 19558
rect 12817 18522 12873 18524
rect 12897 18522 12953 18524
rect 12977 18522 13033 18524
rect 13057 18522 13113 18524
rect 12817 18470 12863 18522
rect 12863 18470 12873 18522
rect 12897 18470 12927 18522
rect 12927 18470 12939 18522
rect 12939 18470 12953 18522
rect 12977 18470 12991 18522
rect 12991 18470 13003 18522
rect 13003 18470 13033 18522
rect 13057 18470 13067 18522
rect 13067 18470 13113 18522
rect 12817 18468 12873 18470
rect 12897 18468 12953 18470
rect 12977 18468 13033 18470
rect 13057 18468 13113 18470
rect 12817 17434 12873 17436
rect 12897 17434 12953 17436
rect 12977 17434 13033 17436
rect 13057 17434 13113 17436
rect 12817 17382 12863 17434
rect 12863 17382 12873 17434
rect 12897 17382 12927 17434
rect 12927 17382 12939 17434
rect 12939 17382 12953 17434
rect 12977 17382 12991 17434
rect 12991 17382 13003 17434
rect 13003 17382 13033 17434
rect 13057 17382 13067 17434
rect 13067 17382 13113 17434
rect 12817 17380 12873 17382
rect 12897 17380 12953 17382
rect 12977 17380 13033 17382
rect 13057 17380 13113 17382
rect 12817 16346 12873 16348
rect 12897 16346 12953 16348
rect 12977 16346 13033 16348
rect 13057 16346 13113 16348
rect 12817 16294 12863 16346
rect 12863 16294 12873 16346
rect 12897 16294 12927 16346
rect 12927 16294 12939 16346
rect 12939 16294 12953 16346
rect 12977 16294 12991 16346
rect 12991 16294 13003 16346
rect 13003 16294 13033 16346
rect 13057 16294 13067 16346
rect 13067 16294 13113 16346
rect 12817 16292 12873 16294
rect 12897 16292 12953 16294
rect 12977 16292 13033 16294
rect 13057 16292 13113 16294
rect 12817 15258 12873 15260
rect 12897 15258 12953 15260
rect 12977 15258 13033 15260
rect 13057 15258 13113 15260
rect 12817 15206 12863 15258
rect 12863 15206 12873 15258
rect 12897 15206 12927 15258
rect 12927 15206 12939 15258
rect 12939 15206 12953 15258
rect 12977 15206 12991 15258
rect 12991 15206 13003 15258
rect 13003 15206 13033 15258
rect 13057 15206 13067 15258
rect 13067 15206 13113 15258
rect 12817 15204 12873 15206
rect 12897 15204 12953 15206
rect 12977 15204 13033 15206
rect 13057 15204 13113 15206
rect 12817 14170 12873 14172
rect 12897 14170 12953 14172
rect 12977 14170 13033 14172
rect 13057 14170 13113 14172
rect 12817 14118 12863 14170
rect 12863 14118 12873 14170
rect 12897 14118 12927 14170
rect 12927 14118 12939 14170
rect 12939 14118 12953 14170
rect 12977 14118 12991 14170
rect 12991 14118 13003 14170
rect 13003 14118 13033 14170
rect 13057 14118 13067 14170
rect 13067 14118 13113 14170
rect 12817 14116 12873 14118
rect 12897 14116 12953 14118
rect 12977 14116 13033 14118
rect 13057 14116 13113 14118
rect 12817 13082 12873 13084
rect 12897 13082 12953 13084
rect 12977 13082 13033 13084
rect 13057 13082 13113 13084
rect 12817 13030 12863 13082
rect 12863 13030 12873 13082
rect 12897 13030 12927 13082
rect 12927 13030 12939 13082
rect 12939 13030 12953 13082
rect 12977 13030 12991 13082
rect 12991 13030 13003 13082
rect 13003 13030 13033 13082
rect 13057 13030 13067 13082
rect 13067 13030 13113 13082
rect 12817 13028 12873 13030
rect 12897 13028 12953 13030
rect 12977 13028 13033 13030
rect 13057 13028 13113 13030
rect 12817 11994 12873 11996
rect 12897 11994 12953 11996
rect 12977 11994 13033 11996
rect 13057 11994 13113 11996
rect 12817 11942 12863 11994
rect 12863 11942 12873 11994
rect 12897 11942 12927 11994
rect 12927 11942 12939 11994
rect 12939 11942 12953 11994
rect 12977 11942 12991 11994
rect 12991 11942 13003 11994
rect 13003 11942 13033 11994
rect 13057 11942 13067 11994
rect 13067 11942 13113 11994
rect 12817 11940 12873 11942
rect 12897 11940 12953 11942
rect 12977 11940 13033 11942
rect 13057 11940 13113 11942
rect 12817 10906 12873 10908
rect 12897 10906 12953 10908
rect 12977 10906 13033 10908
rect 13057 10906 13113 10908
rect 12817 10854 12863 10906
rect 12863 10854 12873 10906
rect 12897 10854 12927 10906
rect 12927 10854 12939 10906
rect 12939 10854 12953 10906
rect 12977 10854 12991 10906
rect 12991 10854 13003 10906
rect 13003 10854 13033 10906
rect 13057 10854 13067 10906
rect 13067 10854 13113 10906
rect 12817 10852 12873 10854
rect 12897 10852 12953 10854
rect 12977 10852 13033 10854
rect 13057 10852 13113 10854
rect 12817 9818 12873 9820
rect 12897 9818 12953 9820
rect 12977 9818 13033 9820
rect 13057 9818 13113 9820
rect 12817 9766 12863 9818
rect 12863 9766 12873 9818
rect 12897 9766 12927 9818
rect 12927 9766 12939 9818
rect 12939 9766 12953 9818
rect 12977 9766 12991 9818
rect 12991 9766 13003 9818
rect 13003 9766 13033 9818
rect 13057 9766 13067 9818
rect 13067 9766 13113 9818
rect 12817 9764 12873 9766
rect 12897 9764 12953 9766
rect 12977 9764 13033 9766
rect 13057 9764 13113 9766
rect 12817 8730 12873 8732
rect 12897 8730 12953 8732
rect 12977 8730 13033 8732
rect 13057 8730 13113 8732
rect 12817 8678 12863 8730
rect 12863 8678 12873 8730
rect 12897 8678 12927 8730
rect 12927 8678 12939 8730
rect 12939 8678 12953 8730
rect 12977 8678 12991 8730
rect 12991 8678 13003 8730
rect 13003 8678 13033 8730
rect 13057 8678 13067 8730
rect 13067 8678 13113 8730
rect 12817 8676 12873 8678
rect 12897 8676 12953 8678
rect 12977 8676 13033 8678
rect 13057 8676 13113 8678
rect 12817 7642 12873 7644
rect 12897 7642 12953 7644
rect 12977 7642 13033 7644
rect 13057 7642 13113 7644
rect 12817 7590 12863 7642
rect 12863 7590 12873 7642
rect 12897 7590 12927 7642
rect 12927 7590 12939 7642
rect 12939 7590 12953 7642
rect 12977 7590 12991 7642
rect 12991 7590 13003 7642
rect 13003 7590 13033 7642
rect 13057 7590 13067 7642
rect 13067 7590 13113 7642
rect 12817 7588 12873 7590
rect 12897 7588 12953 7590
rect 12977 7588 13033 7590
rect 13057 7588 13113 7590
rect 12817 6554 12873 6556
rect 12897 6554 12953 6556
rect 12977 6554 13033 6556
rect 13057 6554 13113 6556
rect 12817 6502 12863 6554
rect 12863 6502 12873 6554
rect 12897 6502 12927 6554
rect 12927 6502 12939 6554
rect 12939 6502 12953 6554
rect 12977 6502 12991 6554
rect 12991 6502 13003 6554
rect 13003 6502 13033 6554
rect 13057 6502 13067 6554
rect 13067 6502 13113 6554
rect 12817 6500 12873 6502
rect 12897 6500 12953 6502
rect 12977 6500 13033 6502
rect 13057 6500 13113 6502
rect 12817 5466 12873 5468
rect 12897 5466 12953 5468
rect 12977 5466 13033 5468
rect 13057 5466 13113 5468
rect 12817 5414 12863 5466
rect 12863 5414 12873 5466
rect 12897 5414 12927 5466
rect 12927 5414 12939 5466
rect 12939 5414 12953 5466
rect 12977 5414 12991 5466
rect 12991 5414 13003 5466
rect 13003 5414 13033 5466
rect 13057 5414 13067 5466
rect 13067 5414 13113 5466
rect 12817 5412 12873 5414
rect 12897 5412 12953 5414
rect 12977 5412 13033 5414
rect 13057 5412 13113 5414
rect 12817 4378 12873 4380
rect 12897 4378 12953 4380
rect 12977 4378 13033 4380
rect 13057 4378 13113 4380
rect 12817 4326 12863 4378
rect 12863 4326 12873 4378
rect 12897 4326 12927 4378
rect 12927 4326 12939 4378
rect 12939 4326 12953 4378
rect 12977 4326 12991 4378
rect 12991 4326 13003 4378
rect 13003 4326 13033 4378
rect 13057 4326 13067 4378
rect 13067 4326 13113 4378
rect 12817 4324 12873 4326
rect 12897 4324 12953 4326
rect 12977 4324 13033 4326
rect 13057 4324 13113 4326
rect 12817 3290 12873 3292
rect 12897 3290 12953 3292
rect 12977 3290 13033 3292
rect 13057 3290 13113 3292
rect 12817 3238 12863 3290
rect 12863 3238 12873 3290
rect 12897 3238 12927 3290
rect 12927 3238 12939 3290
rect 12939 3238 12953 3290
rect 12977 3238 12991 3290
rect 12991 3238 13003 3290
rect 13003 3238 13033 3290
rect 13057 3238 13067 3290
rect 13067 3238 13113 3290
rect 12817 3236 12873 3238
rect 12897 3236 12953 3238
rect 12977 3236 13033 3238
rect 13057 3236 13113 3238
rect 6886 2202 6942 2204
rect 6966 2202 7022 2204
rect 7046 2202 7102 2204
rect 7126 2202 7182 2204
rect 6886 2150 6932 2202
rect 6932 2150 6942 2202
rect 6966 2150 6996 2202
rect 6996 2150 7008 2202
rect 7008 2150 7022 2202
rect 7046 2150 7060 2202
rect 7060 2150 7072 2202
rect 7072 2150 7102 2202
rect 7126 2150 7136 2202
rect 7136 2150 7182 2202
rect 6886 2148 6942 2150
rect 6966 2148 7022 2150
rect 7046 2148 7102 2150
rect 7126 2148 7182 2150
rect 15782 47354 15838 47356
rect 15862 47354 15918 47356
rect 15942 47354 15998 47356
rect 16022 47354 16078 47356
rect 15782 47302 15828 47354
rect 15828 47302 15838 47354
rect 15862 47302 15892 47354
rect 15892 47302 15904 47354
rect 15904 47302 15918 47354
rect 15942 47302 15956 47354
rect 15956 47302 15968 47354
rect 15968 47302 15998 47354
rect 16022 47302 16032 47354
rect 16032 47302 16078 47354
rect 15782 47300 15838 47302
rect 15862 47300 15918 47302
rect 15942 47300 15998 47302
rect 16022 47300 16078 47302
rect 16486 46960 16542 47016
rect 15566 45872 15622 45928
rect 15782 46266 15838 46268
rect 15862 46266 15918 46268
rect 15942 46266 15998 46268
rect 16022 46266 16078 46268
rect 15782 46214 15828 46266
rect 15828 46214 15838 46266
rect 15862 46214 15892 46266
rect 15892 46214 15904 46266
rect 15904 46214 15918 46266
rect 15942 46214 15956 46266
rect 15956 46214 15968 46266
rect 15968 46214 15998 46266
rect 16022 46214 16032 46266
rect 16032 46214 16078 46266
rect 15782 46212 15838 46214
rect 15862 46212 15918 46214
rect 15942 46212 15998 46214
rect 16022 46212 16078 46214
rect 15782 45178 15838 45180
rect 15862 45178 15918 45180
rect 15942 45178 15998 45180
rect 16022 45178 16078 45180
rect 15782 45126 15828 45178
rect 15828 45126 15838 45178
rect 15862 45126 15892 45178
rect 15892 45126 15904 45178
rect 15904 45126 15918 45178
rect 15942 45126 15956 45178
rect 15956 45126 15968 45178
rect 15968 45126 15998 45178
rect 16022 45126 16032 45178
rect 16032 45126 16078 45178
rect 15782 45124 15838 45126
rect 15862 45124 15918 45126
rect 15942 45124 15998 45126
rect 16022 45124 16078 45126
rect 15782 44090 15838 44092
rect 15862 44090 15918 44092
rect 15942 44090 15998 44092
rect 16022 44090 16078 44092
rect 15782 44038 15828 44090
rect 15828 44038 15838 44090
rect 15862 44038 15892 44090
rect 15892 44038 15904 44090
rect 15904 44038 15918 44090
rect 15942 44038 15956 44090
rect 15956 44038 15968 44090
rect 15968 44038 15998 44090
rect 16022 44038 16032 44090
rect 16032 44038 16078 44090
rect 15782 44036 15838 44038
rect 15862 44036 15918 44038
rect 15942 44036 15998 44038
rect 16022 44036 16078 44038
rect 15782 43002 15838 43004
rect 15862 43002 15918 43004
rect 15942 43002 15998 43004
rect 16022 43002 16078 43004
rect 15782 42950 15828 43002
rect 15828 42950 15838 43002
rect 15862 42950 15892 43002
rect 15892 42950 15904 43002
rect 15904 42950 15918 43002
rect 15942 42950 15956 43002
rect 15956 42950 15968 43002
rect 15968 42950 15998 43002
rect 16022 42950 16032 43002
rect 16032 42950 16078 43002
rect 15782 42948 15838 42950
rect 15862 42948 15918 42950
rect 15942 42948 15998 42950
rect 16022 42948 16078 42950
rect 15782 41914 15838 41916
rect 15862 41914 15918 41916
rect 15942 41914 15998 41916
rect 16022 41914 16078 41916
rect 15782 41862 15828 41914
rect 15828 41862 15838 41914
rect 15862 41862 15892 41914
rect 15892 41862 15904 41914
rect 15904 41862 15918 41914
rect 15942 41862 15956 41914
rect 15956 41862 15968 41914
rect 15968 41862 15998 41914
rect 16022 41862 16032 41914
rect 16032 41862 16078 41914
rect 15782 41860 15838 41862
rect 15862 41860 15918 41862
rect 15942 41860 15998 41862
rect 16022 41860 16078 41862
rect 15782 40826 15838 40828
rect 15862 40826 15918 40828
rect 15942 40826 15998 40828
rect 16022 40826 16078 40828
rect 15782 40774 15828 40826
rect 15828 40774 15838 40826
rect 15862 40774 15892 40826
rect 15892 40774 15904 40826
rect 15904 40774 15918 40826
rect 15942 40774 15956 40826
rect 15956 40774 15968 40826
rect 15968 40774 15998 40826
rect 16022 40774 16032 40826
rect 16032 40774 16078 40826
rect 15782 40772 15838 40774
rect 15862 40772 15918 40774
rect 15942 40772 15998 40774
rect 16022 40772 16078 40774
rect 15782 39738 15838 39740
rect 15862 39738 15918 39740
rect 15942 39738 15998 39740
rect 16022 39738 16078 39740
rect 15782 39686 15828 39738
rect 15828 39686 15838 39738
rect 15862 39686 15892 39738
rect 15892 39686 15904 39738
rect 15904 39686 15918 39738
rect 15942 39686 15956 39738
rect 15956 39686 15968 39738
rect 15968 39686 15998 39738
rect 16022 39686 16032 39738
rect 16032 39686 16078 39738
rect 15782 39684 15838 39686
rect 15862 39684 15918 39686
rect 15942 39684 15998 39686
rect 16022 39684 16078 39686
rect 15782 38650 15838 38652
rect 15862 38650 15918 38652
rect 15942 38650 15998 38652
rect 16022 38650 16078 38652
rect 15782 38598 15828 38650
rect 15828 38598 15838 38650
rect 15862 38598 15892 38650
rect 15892 38598 15904 38650
rect 15904 38598 15918 38650
rect 15942 38598 15956 38650
rect 15956 38598 15968 38650
rect 15968 38598 15998 38650
rect 16022 38598 16032 38650
rect 16032 38598 16078 38650
rect 15782 38596 15838 38598
rect 15862 38596 15918 38598
rect 15942 38596 15998 38598
rect 16022 38596 16078 38598
rect 15782 37562 15838 37564
rect 15862 37562 15918 37564
rect 15942 37562 15998 37564
rect 16022 37562 16078 37564
rect 15782 37510 15828 37562
rect 15828 37510 15838 37562
rect 15862 37510 15892 37562
rect 15892 37510 15904 37562
rect 15904 37510 15918 37562
rect 15942 37510 15956 37562
rect 15956 37510 15968 37562
rect 15968 37510 15998 37562
rect 16022 37510 16032 37562
rect 16032 37510 16078 37562
rect 15782 37508 15838 37510
rect 15862 37508 15918 37510
rect 15942 37508 15998 37510
rect 16022 37508 16078 37510
rect 15782 36474 15838 36476
rect 15862 36474 15918 36476
rect 15942 36474 15998 36476
rect 16022 36474 16078 36476
rect 15782 36422 15828 36474
rect 15828 36422 15838 36474
rect 15862 36422 15892 36474
rect 15892 36422 15904 36474
rect 15904 36422 15918 36474
rect 15942 36422 15956 36474
rect 15956 36422 15968 36474
rect 15968 36422 15998 36474
rect 16022 36422 16032 36474
rect 16032 36422 16078 36474
rect 15782 36420 15838 36422
rect 15862 36420 15918 36422
rect 15942 36420 15998 36422
rect 16022 36420 16078 36422
rect 15782 35386 15838 35388
rect 15862 35386 15918 35388
rect 15942 35386 15998 35388
rect 16022 35386 16078 35388
rect 15782 35334 15828 35386
rect 15828 35334 15838 35386
rect 15862 35334 15892 35386
rect 15892 35334 15904 35386
rect 15904 35334 15918 35386
rect 15942 35334 15956 35386
rect 15956 35334 15968 35386
rect 15968 35334 15998 35386
rect 16022 35334 16032 35386
rect 16032 35334 16078 35386
rect 15782 35332 15838 35334
rect 15862 35332 15918 35334
rect 15942 35332 15998 35334
rect 16022 35332 16078 35334
rect 15750 34584 15806 34640
rect 15658 34448 15714 34504
rect 15782 34298 15838 34300
rect 15862 34298 15918 34300
rect 15942 34298 15998 34300
rect 16022 34298 16078 34300
rect 15782 34246 15828 34298
rect 15828 34246 15838 34298
rect 15862 34246 15892 34298
rect 15892 34246 15904 34298
rect 15904 34246 15918 34298
rect 15942 34246 15956 34298
rect 15956 34246 15968 34298
rect 15968 34246 15998 34298
rect 16022 34246 16032 34298
rect 16032 34246 16078 34298
rect 15782 34244 15838 34246
rect 15862 34244 15918 34246
rect 15942 34244 15998 34246
rect 16022 34244 16078 34246
rect 15566 33496 15622 33552
rect 15782 33210 15838 33212
rect 15862 33210 15918 33212
rect 15942 33210 15998 33212
rect 16022 33210 16078 33212
rect 15782 33158 15828 33210
rect 15828 33158 15838 33210
rect 15862 33158 15892 33210
rect 15892 33158 15904 33210
rect 15904 33158 15918 33210
rect 15942 33158 15956 33210
rect 15956 33158 15968 33210
rect 15968 33158 15998 33210
rect 16022 33158 16032 33210
rect 16032 33158 16078 33210
rect 15782 33156 15838 33158
rect 15862 33156 15918 33158
rect 15942 33156 15998 33158
rect 16022 33156 16078 33158
rect 15782 32122 15838 32124
rect 15862 32122 15918 32124
rect 15942 32122 15998 32124
rect 16022 32122 16078 32124
rect 15782 32070 15828 32122
rect 15828 32070 15838 32122
rect 15862 32070 15892 32122
rect 15892 32070 15904 32122
rect 15904 32070 15918 32122
rect 15942 32070 15956 32122
rect 15956 32070 15968 32122
rect 15968 32070 15998 32122
rect 16022 32070 16032 32122
rect 16032 32070 16078 32122
rect 15782 32068 15838 32070
rect 15862 32068 15918 32070
rect 15942 32068 15998 32070
rect 16022 32068 16078 32070
rect 15782 31034 15838 31036
rect 15862 31034 15918 31036
rect 15942 31034 15998 31036
rect 16022 31034 16078 31036
rect 15782 30982 15828 31034
rect 15828 30982 15838 31034
rect 15862 30982 15892 31034
rect 15892 30982 15904 31034
rect 15904 30982 15918 31034
rect 15942 30982 15956 31034
rect 15956 30982 15968 31034
rect 15968 30982 15998 31034
rect 16022 30982 16032 31034
rect 16032 30982 16078 31034
rect 15782 30980 15838 30982
rect 15862 30980 15918 30982
rect 15942 30980 15998 30982
rect 16022 30980 16078 30982
rect 15782 29946 15838 29948
rect 15862 29946 15918 29948
rect 15942 29946 15998 29948
rect 16022 29946 16078 29948
rect 15782 29894 15828 29946
rect 15828 29894 15838 29946
rect 15862 29894 15892 29946
rect 15892 29894 15904 29946
rect 15904 29894 15918 29946
rect 15942 29894 15956 29946
rect 15956 29894 15968 29946
rect 15968 29894 15998 29946
rect 16022 29894 16032 29946
rect 16032 29894 16078 29946
rect 15782 29892 15838 29894
rect 15862 29892 15918 29894
rect 15942 29892 15998 29894
rect 16022 29892 16078 29894
rect 15782 28858 15838 28860
rect 15862 28858 15918 28860
rect 15942 28858 15998 28860
rect 16022 28858 16078 28860
rect 15782 28806 15828 28858
rect 15828 28806 15838 28858
rect 15862 28806 15892 28858
rect 15892 28806 15904 28858
rect 15904 28806 15918 28858
rect 15942 28806 15956 28858
rect 15956 28806 15968 28858
rect 15968 28806 15998 28858
rect 16022 28806 16032 28858
rect 16032 28806 16078 28858
rect 15782 28804 15838 28806
rect 15862 28804 15918 28806
rect 15942 28804 15998 28806
rect 16022 28804 16078 28806
rect 16578 33224 16634 33280
rect 16946 34604 17002 34640
rect 16946 34584 16948 34604
rect 16948 34584 17000 34604
rect 17000 34584 17002 34604
rect 18142 40704 18198 40760
rect 17590 33496 17646 33552
rect 15782 27770 15838 27772
rect 15862 27770 15918 27772
rect 15942 27770 15998 27772
rect 16022 27770 16078 27772
rect 15782 27718 15828 27770
rect 15828 27718 15838 27770
rect 15862 27718 15892 27770
rect 15892 27718 15904 27770
rect 15904 27718 15918 27770
rect 15942 27718 15956 27770
rect 15956 27718 15968 27770
rect 15968 27718 15998 27770
rect 16022 27718 16032 27770
rect 16032 27718 16078 27770
rect 15782 27716 15838 27718
rect 15862 27716 15918 27718
rect 15942 27716 15998 27718
rect 16022 27716 16078 27718
rect 15782 26682 15838 26684
rect 15862 26682 15918 26684
rect 15942 26682 15998 26684
rect 16022 26682 16078 26684
rect 15782 26630 15828 26682
rect 15828 26630 15838 26682
rect 15862 26630 15892 26682
rect 15892 26630 15904 26682
rect 15904 26630 15918 26682
rect 15942 26630 15956 26682
rect 15956 26630 15968 26682
rect 15968 26630 15998 26682
rect 16022 26630 16032 26682
rect 16032 26630 16078 26682
rect 15782 26628 15838 26630
rect 15862 26628 15918 26630
rect 15942 26628 15998 26630
rect 16022 26628 16078 26630
rect 15782 25594 15838 25596
rect 15862 25594 15918 25596
rect 15942 25594 15998 25596
rect 16022 25594 16078 25596
rect 15782 25542 15828 25594
rect 15828 25542 15838 25594
rect 15862 25542 15892 25594
rect 15892 25542 15904 25594
rect 15904 25542 15918 25594
rect 15942 25542 15956 25594
rect 15956 25542 15968 25594
rect 15968 25542 15998 25594
rect 16022 25542 16032 25594
rect 16032 25542 16078 25594
rect 15782 25540 15838 25542
rect 15862 25540 15918 25542
rect 15942 25540 15998 25542
rect 16022 25540 16078 25542
rect 15782 24506 15838 24508
rect 15862 24506 15918 24508
rect 15942 24506 15998 24508
rect 16022 24506 16078 24508
rect 15782 24454 15828 24506
rect 15828 24454 15838 24506
rect 15862 24454 15892 24506
rect 15892 24454 15904 24506
rect 15904 24454 15918 24506
rect 15942 24454 15956 24506
rect 15956 24454 15968 24506
rect 15968 24454 15998 24506
rect 16022 24454 16032 24506
rect 16032 24454 16078 24506
rect 15782 24452 15838 24454
rect 15862 24452 15918 24454
rect 15942 24452 15998 24454
rect 16022 24452 16078 24454
rect 15782 23418 15838 23420
rect 15862 23418 15918 23420
rect 15942 23418 15998 23420
rect 16022 23418 16078 23420
rect 15782 23366 15828 23418
rect 15828 23366 15838 23418
rect 15862 23366 15892 23418
rect 15892 23366 15904 23418
rect 15904 23366 15918 23418
rect 15942 23366 15956 23418
rect 15956 23366 15968 23418
rect 15968 23366 15998 23418
rect 16022 23366 16032 23418
rect 16032 23366 16078 23418
rect 15782 23364 15838 23366
rect 15862 23364 15918 23366
rect 15942 23364 15998 23366
rect 16022 23364 16078 23366
rect 15782 22330 15838 22332
rect 15862 22330 15918 22332
rect 15942 22330 15998 22332
rect 16022 22330 16078 22332
rect 15782 22278 15828 22330
rect 15828 22278 15838 22330
rect 15862 22278 15892 22330
rect 15892 22278 15904 22330
rect 15904 22278 15918 22330
rect 15942 22278 15956 22330
rect 15956 22278 15968 22330
rect 15968 22278 15998 22330
rect 16022 22278 16032 22330
rect 16032 22278 16078 22330
rect 15782 22276 15838 22278
rect 15862 22276 15918 22278
rect 15942 22276 15998 22278
rect 16022 22276 16078 22278
rect 15782 21242 15838 21244
rect 15862 21242 15918 21244
rect 15942 21242 15998 21244
rect 16022 21242 16078 21244
rect 15782 21190 15828 21242
rect 15828 21190 15838 21242
rect 15862 21190 15892 21242
rect 15892 21190 15904 21242
rect 15904 21190 15918 21242
rect 15942 21190 15956 21242
rect 15956 21190 15968 21242
rect 15968 21190 15998 21242
rect 16022 21190 16032 21242
rect 16032 21190 16078 21242
rect 15782 21188 15838 21190
rect 15862 21188 15918 21190
rect 15942 21188 15998 21190
rect 16022 21188 16078 21190
rect 15782 20154 15838 20156
rect 15862 20154 15918 20156
rect 15942 20154 15998 20156
rect 16022 20154 16078 20156
rect 15782 20102 15828 20154
rect 15828 20102 15838 20154
rect 15862 20102 15892 20154
rect 15892 20102 15904 20154
rect 15904 20102 15918 20154
rect 15942 20102 15956 20154
rect 15956 20102 15968 20154
rect 15968 20102 15998 20154
rect 16022 20102 16032 20154
rect 16032 20102 16078 20154
rect 15782 20100 15838 20102
rect 15862 20100 15918 20102
rect 15942 20100 15998 20102
rect 16022 20100 16078 20102
rect 15782 19066 15838 19068
rect 15862 19066 15918 19068
rect 15942 19066 15998 19068
rect 16022 19066 16078 19068
rect 15782 19014 15828 19066
rect 15828 19014 15838 19066
rect 15862 19014 15892 19066
rect 15892 19014 15904 19066
rect 15904 19014 15918 19066
rect 15942 19014 15956 19066
rect 15956 19014 15968 19066
rect 15968 19014 15998 19066
rect 16022 19014 16032 19066
rect 16032 19014 16078 19066
rect 15782 19012 15838 19014
rect 15862 19012 15918 19014
rect 15942 19012 15998 19014
rect 16022 19012 16078 19014
rect 15782 17978 15838 17980
rect 15862 17978 15918 17980
rect 15942 17978 15998 17980
rect 16022 17978 16078 17980
rect 15782 17926 15828 17978
rect 15828 17926 15838 17978
rect 15862 17926 15892 17978
rect 15892 17926 15904 17978
rect 15904 17926 15918 17978
rect 15942 17926 15956 17978
rect 15956 17926 15968 17978
rect 15968 17926 15998 17978
rect 16022 17926 16032 17978
rect 16032 17926 16078 17978
rect 15782 17924 15838 17926
rect 15862 17924 15918 17926
rect 15942 17924 15998 17926
rect 16022 17924 16078 17926
rect 15782 16890 15838 16892
rect 15862 16890 15918 16892
rect 15942 16890 15998 16892
rect 16022 16890 16078 16892
rect 15782 16838 15828 16890
rect 15828 16838 15838 16890
rect 15862 16838 15892 16890
rect 15892 16838 15904 16890
rect 15904 16838 15918 16890
rect 15942 16838 15956 16890
rect 15956 16838 15968 16890
rect 15968 16838 15998 16890
rect 16022 16838 16032 16890
rect 16032 16838 16078 16890
rect 15782 16836 15838 16838
rect 15862 16836 15918 16838
rect 15942 16836 15998 16838
rect 16022 16836 16078 16838
rect 15782 15802 15838 15804
rect 15862 15802 15918 15804
rect 15942 15802 15998 15804
rect 16022 15802 16078 15804
rect 15782 15750 15828 15802
rect 15828 15750 15838 15802
rect 15862 15750 15892 15802
rect 15892 15750 15904 15802
rect 15904 15750 15918 15802
rect 15942 15750 15956 15802
rect 15956 15750 15968 15802
rect 15968 15750 15998 15802
rect 16022 15750 16032 15802
rect 16032 15750 16078 15802
rect 15782 15748 15838 15750
rect 15862 15748 15918 15750
rect 15942 15748 15998 15750
rect 16022 15748 16078 15750
rect 15782 14714 15838 14716
rect 15862 14714 15918 14716
rect 15942 14714 15998 14716
rect 16022 14714 16078 14716
rect 15782 14662 15828 14714
rect 15828 14662 15838 14714
rect 15862 14662 15892 14714
rect 15892 14662 15904 14714
rect 15904 14662 15918 14714
rect 15942 14662 15956 14714
rect 15956 14662 15968 14714
rect 15968 14662 15998 14714
rect 16022 14662 16032 14714
rect 16032 14662 16078 14714
rect 15782 14660 15838 14662
rect 15862 14660 15918 14662
rect 15942 14660 15998 14662
rect 16022 14660 16078 14662
rect 15782 13626 15838 13628
rect 15862 13626 15918 13628
rect 15942 13626 15998 13628
rect 16022 13626 16078 13628
rect 15782 13574 15828 13626
rect 15828 13574 15838 13626
rect 15862 13574 15892 13626
rect 15892 13574 15904 13626
rect 15904 13574 15918 13626
rect 15942 13574 15956 13626
rect 15956 13574 15968 13626
rect 15968 13574 15998 13626
rect 16022 13574 16032 13626
rect 16032 13574 16078 13626
rect 15782 13572 15838 13574
rect 15862 13572 15918 13574
rect 15942 13572 15998 13574
rect 16022 13572 16078 13574
rect 15782 12538 15838 12540
rect 15862 12538 15918 12540
rect 15942 12538 15998 12540
rect 16022 12538 16078 12540
rect 15782 12486 15828 12538
rect 15828 12486 15838 12538
rect 15862 12486 15892 12538
rect 15892 12486 15904 12538
rect 15904 12486 15918 12538
rect 15942 12486 15956 12538
rect 15956 12486 15968 12538
rect 15968 12486 15998 12538
rect 16022 12486 16032 12538
rect 16032 12486 16078 12538
rect 15782 12484 15838 12486
rect 15862 12484 15918 12486
rect 15942 12484 15998 12486
rect 16022 12484 16078 12486
rect 15782 11450 15838 11452
rect 15862 11450 15918 11452
rect 15942 11450 15998 11452
rect 16022 11450 16078 11452
rect 15782 11398 15828 11450
rect 15828 11398 15838 11450
rect 15862 11398 15892 11450
rect 15892 11398 15904 11450
rect 15904 11398 15918 11450
rect 15942 11398 15956 11450
rect 15956 11398 15968 11450
rect 15968 11398 15998 11450
rect 16022 11398 16032 11450
rect 16032 11398 16078 11450
rect 15782 11396 15838 11398
rect 15862 11396 15918 11398
rect 15942 11396 15998 11398
rect 16022 11396 16078 11398
rect 15782 10362 15838 10364
rect 15862 10362 15918 10364
rect 15942 10362 15998 10364
rect 16022 10362 16078 10364
rect 15782 10310 15828 10362
rect 15828 10310 15838 10362
rect 15862 10310 15892 10362
rect 15892 10310 15904 10362
rect 15904 10310 15918 10362
rect 15942 10310 15956 10362
rect 15956 10310 15968 10362
rect 15968 10310 15998 10362
rect 16022 10310 16032 10362
rect 16032 10310 16078 10362
rect 15782 10308 15838 10310
rect 15862 10308 15918 10310
rect 15942 10308 15998 10310
rect 16022 10308 16078 10310
rect 15782 9274 15838 9276
rect 15862 9274 15918 9276
rect 15942 9274 15998 9276
rect 16022 9274 16078 9276
rect 15782 9222 15828 9274
rect 15828 9222 15838 9274
rect 15862 9222 15892 9274
rect 15892 9222 15904 9274
rect 15904 9222 15918 9274
rect 15942 9222 15956 9274
rect 15956 9222 15968 9274
rect 15968 9222 15998 9274
rect 16022 9222 16032 9274
rect 16032 9222 16078 9274
rect 15782 9220 15838 9222
rect 15862 9220 15918 9222
rect 15942 9220 15998 9222
rect 16022 9220 16078 9222
rect 15782 8186 15838 8188
rect 15862 8186 15918 8188
rect 15942 8186 15998 8188
rect 16022 8186 16078 8188
rect 15782 8134 15828 8186
rect 15828 8134 15838 8186
rect 15862 8134 15892 8186
rect 15892 8134 15904 8186
rect 15904 8134 15918 8186
rect 15942 8134 15956 8186
rect 15956 8134 15968 8186
rect 15968 8134 15998 8186
rect 16022 8134 16032 8186
rect 16032 8134 16078 8186
rect 15782 8132 15838 8134
rect 15862 8132 15918 8134
rect 15942 8132 15998 8134
rect 16022 8132 16078 8134
rect 15782 7098 15838 7100
rect 15862 7098 15918 7100
rect 15942 7098 15998 7100
rect 16022 7098 16078 7100
rect 15782 7046 15828 7098
rect 15828 7046 15838 7098
rect 15862 7046 15892 7098
rect 15892 7046 15904 7098
rect 15904 7046 15918 7098
rect 15942 7046 15956 7098
rect 15956 7046 15968 7098
rect 15968 7046 15998 7098
rect 16022 7046 16032 7098
rect 16032 7046 16078 7098
rect 15782 7044 15838 7046
rect 15862 7044 15918 7046
rect 15942 7044 15998 7046
rect 16022 7044 16078 7046
rect 15782 6010 15838 6012
rect 15862 6010 15918 6012
rect 15942 6010 15998 6012
rect 16022 6010 16078 6012
rect 15782 5958 15828 6010
rect 15828 5958 15838 6010
rect 15862 5958 15892 6010
rect 15892 5958 15904 6010
rect 15904 5958 15918 6010
rect 15942 5958 15956 6010
rect 15956 5958 15968 6010
rect 15968 5958 15998 6010
rect 16022 5958 16032 6010
rect 16032 5958 16078 6010
rect 15782 5956 15838 5958
rect 15862 5956 15918 5958
rect 15942 5956 15998 5958
rect 16022 5956 16078 5958
rect 15782 4922 15838 4924
rect 15862 4922 15918 4924
rect 15942 4922 15998 4924
rect 16022 4922 16078 4924
rect 15782 4870 15828 4922
rect 15828 4870 15838 4922
rect 15862 4870 15892 4922
rect 15892 4870 15904 4922
rect 15904 4870 15918 4922
rect 15942 4870 15956 4922
rect 15956 4870 15968 4922
rect 15968 4870 15998 4922
rect 16022 4870 16032 4922
rect 16032 4870 16078 4922
rect 15782 4868 15838 4870
rect 15862 4868 15918 4870
rect 15942 4868 15998 4870
rect 16022 4868 16078 4870
rect 15782 3834 15838 3836
rect 15862 3834 15918 3836
rect 15942 3834 15998 3836
rect 16022 3834 16078 3836
rect 15782 3782 15828 3834
rect 15828 3782 15838 3834
rect 15862 3782 15892 3834
rect 15892 3782 15904 3834
rect 15904 3782 15918 3834
rect 15942 3782 15956 3834
rect 15956 3782 15968 3834
rect 15968 3782 15998 3834
rect 16022 3782 16032 3834
rect 16032 3782 16078 3834
rect 15782 3780 15838 3782
rect 15862 3780 15918 3782
rect 15942 3780 15998 3782
rect 16022 3780 16078 3782
rect 18142 28192 18198 28248
rect 18142 21972 18144 21992
rect 18144 21972 18196 21992
rect 18196 21972 18198 21992
rect 18142 21936 18198 21972
rect 18142 15700 18198 15736
rect 18142 15680 18144 15700
rect 18144 15680 18196 15700
rect 18196 15680 18198 15700
rect 18050 9444 18106 9480
rect 18050 9424 18052 9444
rect 18052 9424 18104 9444
rect 18104 9424 18106 9444
rect 18050 3168 18106 3224
rect 15782 2746 15838 2748
rect 15862 2746 15918 2748
rect 15942 2746 15998 2748
rect 16022 2746 16078 2748
rect 15782 2694 15828 2746
rect 15828 2694 15838 2746
rect 15862 2694 15892 2746
rect 15892 2694 15904 2746
rect 15904 2694 15918 2746
rect 15942 2694 15956 2746
rect 15956 2694 15968 2746
rect 15968 2694 15998 2746
rect 16022 2694 16032 2746
rect 16032 2694 16078 2746
rect 15782 2692 15838 2694
rect 15862 2692 15918 2694
rect 15942 2692 15998 2694
rect 16022 2692 16078 2694
rect 12817 2202 12873 2204
rect 12897 2202 12953 2204
rect 12977 2202 13033 2204
rect 13057 2202 13113 2204
rect 12817 2150 12863 2202
rect 12863 2150 12873 2202
rect 12897 2150 12927 2202
rect 12927 2150 12939 2202
rect 12939 2150 12953 2202
rect 12977 2150 12991 2202
rect 12991 2150 13003 2202
rect 13003 2150 13033 2202
rect 13057 2150 13067 2202
rect 13067 2150 13113 2202
rect 12817 2148 12873 2150
rect 12897 2148 12953 2150
rect 12977 2148 13033 2150
rect 13057 2148 13113 2150
<< metal3 >>
rect 3909 47360 4229 47361
rect 0 47290 800 47320
rect 3909 47296 3917 47360
rect 3981 47296 3997 47360
rect 4061 47296 4077 47360
rect 4141 47296 4157 47360
rect 4221 47296 4229 47360
rect 3909 47295 4229 47296
rect 9840 47360 10160 47361
rect 9840 47296 9848 47360
rect 9912 47296 9928 47360
rect 9992 47296 10008 47360
rect 10072 47296 10088 47360
rect 10152 47296 10160 47360
rect 9840 47295 10160 47296
rect 15770 47360 16090 47361
rect 15770 47296 15778 47360
rect 15842 47296 15858 47360
rect 15922 47296 15938 47360
rect 16002 47296 16018 47360
rect 16082 47296 16090 47360
rect 15770 47295 16090 47296
rect 1485 47290 1551 47293
rect 0 47288 1551 47290
rect 0 47232 1490 47288
rect 1546 47232 1551 47288
rect 0 47230 1551 47232
rect 0 47200 800 47230
rect 1485 47227 1551 47230
rect 16481 47018 16547 47021
rect 19200 47018 20000 47048
rect 16481 47016 20000 47018
rect 16481 46960 16486 47016
rect 16542 46960 20000 47016
rect 16481 46958 20000 46960
rect 16481 46955 16547 46958
rect 19200 46928 20000 46958
rect 6874 46816 7194 46817
rect 6874 46752 6882 46816
rect 6946 46752 6962 46816
rect 7026 46752 7042 46816
rect 7106 46752 7122 46816
rect 7186 46752 7194 46816
rect 6874 46751 7194 46752
rect 12805 46816 13125 46817
rect 12805 46752 12813 46816
rect 12877 46752 12893 46816
rect 12957 46752 12973 46816
rect 13037 46752 13053 46816
rect 13117 46752 13125 46816
rect 12805 46751 13125 46752
rect 3909 46272 4229 46273
rect 3909 46208 3917 46272
rect 3981 46208 3997 46272
rect 4061 46208 4077 46272
rect 4141 46208 4157 46272
rect 4221 46208 4229 46272
rect 3909 46207 4229 46208
rect 9840 46272 10160 46273
rect 9840 46208 9848 46272
rect 9912 46208 9928 46272
rect 9992 46208 10008 46272
rect 10072 46208 10088 46272
rect 10152 46208 10160 46272
rect 9840 46207 10160 46208
rect 15770 46272 16090 46273
rect 15770 46208 15778 46272
rect 15842 46208 15858 46272
rect 15922 46208 15938 46272
rect 16002 46208 16018 46272
rect 16082 46208 16090 46272
rect 15770 46207 16090 46208
rect 15561 45932 15627 45933
rect 15510 45930 15516 45932
rect 15470 45870 15516 45930
rect 15580 45928 15627 45932
rect 15622 45872 15627 45928
rect 15510 45868 15516 45870
rect 15580 45868 15627 45872
rect 15561 45867 15627 45868
rect 6874 45728 7194 45729
rect 6874 45664 6882 45728
rect 6946 45664 6962 45728
rect 7026 45664 7042 45728
rect 7106 45664 7122 45728
rect 7186 45664 7194 45728
rect 6874 45663 7194 45664
rect 12805 45728 13125 45729
rect 12805 45664 12813 45728
rect 12877 45664 12893 45728
rect 12957 45664 12973 45728
rect 13037 45664 13053 45728
rect 13117 45664 13125 45728
rect 12805 45663 13125 45664
rect 3909 45184 4229 45185
rect 3909 45120 3917 45184
rect 3981 45120 3997 45184
rect 4061 45120 4077 45184
rect 4141 45120 4157 45184
rect 4221 45120 4229 45184
rect 3909 45119 4229 45120
rect 9840 45184 10160 45185
rect 9840 45120 9848 45184
rect 9912 45120 9928 45184
rect 9992 45120 10008 45184
rect 10072 45120 10088 45184
rect 10152 45120 10160 45184
rect 9840 45119 10160 45120
rect 15770 45184 16090 45185
rect 15770 45120 15778 45184
rect 15842 45120 15858 45184
rect 15922 45120 15938 45184
rect 16002 45120 16018 45184
rect 16082 45120 16090 45184
rect 15770 45119 16090 45120
rect 6874 44640 7194 44641
rect 6874 44576 6882 44640
rect 6946 44576 6962 44640
rect 7026 44576 7042 44640
rect 7106 44576 7122 44640
rect 7186 44576 7194 44640
rect 6874 44575 7194 44576
rect 12805 44640 13125 44641
rect 12805 44576 12813 44640
rect 12877 44576 12893 44640
rect 12957 44576 12973 44640
rect 13037 44576 13053 44640
rect 13117 44576 13125 44640
rect 12805 44575 13125 44576
rect 3909 44096 4229 44097
rect 3909 44032 3917 44096
rect 3981 44032 3997 44096
rect 4061 44032 4077 44096
rect 4141 44032 4157 44096
rect 4221 44032 4229 44096
rect 3909 44031 4229 44032
rect 9840 44096 10160 44097
rect 9840 44032 9848 44096
rect 9912 44032 9928 44096
rect 9992 44032 10008 44096
rect 10072 44032 10088 44096
rect 10152 44032 10160 44096
rect 9840 44031 10160 44032
rect 15770 44096 16090 44097
rect 15770 44032 15778 44096
rect 15842 44032 15858 44096
rect 15922 44032 15938 44096
rect 16002 44032 16018 44096
rect 16082 44032 16090 44096
rect 15770 44031 16090 44032
rect 6874 43552 7194 43553
rect 6874 43488 6882 43552
rect 6946 43488 6962 43552
rect 7026 43488 7042 43552
rect 7106 43488 7122 43552
rect 7186 43488 7194 43552
rect 6874 43487 7194 43488
rect 12805 43552 13125 43553
rect 12805 43488 12813 43552
rect 12877 43488 12893 43552
rect 12957 43488 12973 43552
rect 13037 43488 13053 43552
rect 13117 43488 13125 43552
rect 12805 43487 13125 43488
rect 3909 43008 4229 43009
rect 3909 42944 3917 43008
rect 3981 42944 3997 43008
rect 4061 42944 4077 43008
rect 4141 42944 4157 43008
rect 4221 42944 4229 43008
rect 3909 42943 4229 42944
rect 9840 43008 10160 43009
rect 9840 42944 9848 43008
rect 9912 42944 9928 43008
rect 9992 42944 10008 43008
rect 10072 42944 10088 43008
rect 10152 42944 10160 43008
rect 9840 42943 10160 42944
rect 15770 43008 16090 43009
rect 15770 42944 15778 43008
rect 15842 42944 15858 43008
rect 15922 42944 15938 43008
rect 16002 42944 16018 43008
rect 16082 42944 16090 43008
rect 15770 42943 16090 42944
rect 6874 42464 7194 42465
rect 6874 42400 6882 42464
rect 6946 42400 6962 42464
rect 7026 42400 7042 42464
rect 7106 42400 7122 42464
rect 7186 42400 7194 42464
rect 6874 42399 7194 42400
rect 12805 42464 13125 42465
rect 12805 42400 12813 42464
rect 12877 42400 12893 42464
rect 12957 42400 12973 42464
rect 13037 42400 13053 42464
rect 13117 42400 13125 42464
rect 12805 42399 13125 42400
rect 3909 41920 4229 41921
rect 3909 41856 3917 41920
rect 3981 41856 3997 41920
rect 4061 41856 4077 41920
rect 4141 41856 4157 41920
rect 4221 41856 4229 41920
rect 3909 41855 4229 41856
rect 9840 41920 10160 41921
rect 9840 41856 9848 41920
rect 9912 41856 9928 41920
rect 9992 41856 10008 41920
rect 10072 41856 10088 41920
rect 10152 41856 10160 41920
rect 9840 41855 10160 41856
rect 15770 41920 16090 41921
rect 15770 41856 15778 41920
rect 15842 41856 15858 41920
rect 15922 41856 15938 41920
rect 16002 41856 16018 41920
rect 16082 41856 16090 41920
rect 15770 41855 16090 41856
rect 0 41714 800 41744
rect 1485 41714 1551 41717
rect 0 41712 1551 41714
rect 0 41656 1490 41712
rect 1546 41656 1551 41712
rect 0 41654 1551 41656
rect 0 41624 800 41654
rect 1485 41651 1551 41654
rect 6874 41376 7194 41377
rect 6874 41312 6882 41376
rect 6946 41312 6962 41376
rect 7026 41312 7042 41376
rect 7106 41312 7122 41376
rect 7186 41312 7194 41376
rect 6874 41311 7194 41312
rect 12805 41376 13125 41377
rect 12805 41312 12813 41376
rect 12877 41312 12893 41376
rect 12957 41312 12973 41376
rect 13037 41312 13053 41376
rect 13117 41312 13125 41376
rect 12805 41311 13125 41312
rect 3909 40832 4229 40833
rect 3909 40768 3917 40832
rect 3981 40768 3997 40832
rect 4061 40768 4077 40832
rect 4141 40768 4157 40832
rect 4221 40768 4229 40832
rect 3909 40767 4229 40768
rect 9840 40832 10160 40833
rect 9840 40768 9848 40832
rect 9912 40768 9928 40832
rect 9992 40768 10008 40832
rect 10072 40768 10088 40832
rect 10152 40768 10160 40832
rect 9840 40767 10160 40768
rect 15770 40832 16090 40833
rect 15770 40768 15778 40832
rect 15842 40768 15858 40832
rect 15922 40768 15938 40832
rect 16002 40768 16018 40832
rect 16082 40768 16090 40832
rect 15770 40767 16090 40768
rect 18137 40762 18203 40765
rect 19200 40762 20000 40792
rect 18137 40760 20000 40762
rect 18137 40704 18142 40760
rect 18198 40704 20000 40760
rect 18137 40702 20000 40704
rect 18137 40699 18203 40702
rect 19200 40672 20000 40702
rect 6874 40288 7194 40289
rect 6874 40224 6882 40288
rect 6946 40224 6962 40288
rect 7026 40224 7042 40288
rect 7106 40224 7122 40288
rect 7186 40224 7194 40288
rect 6874 40223 7194 40224
rect 12805 40288 13125 40289
rect 12805 40224 12813 40288
rect 12877 40224 12893 40288
rect 12957 40224 12973 40288
rect 13037 40224 13053 40288
rect 13117 40224 13125 40288
rect 12805 40223 13125 40224
rect 3909 39744 4229 39745
rect 3909 39680 3917 39744
rect 3981 39680 3997 39744
rect 4061 39680 4077 39744
rect 4141 39680 4157 39744
rect 4221 39680 4229 39744
rect 3909 39679 4229 39680
rect 9840 39744 10160 39745
rect 9840 39680 9848 39744
rect 9912 39680 9928 39744
rect 9992 39680 10008 39744
rect 10072 39680 10088 39744
rect 10152 39680 10160 39744
rect 9840 39679 10160 39680
rect 15770 39744 16090 39745
rect 15770 39680 15778 39744
rect 15842 39680 15858 39744
rect 15922 39680 15938 39744
rect 16002 39680 16018 39744
rect 16082 39680 16090 39744
rect 15770 39679 16090 39680
rect 6874 39200 7194 39201
rect 6874 39136 6882 39200
rect 6946 39136 6962 39200
rect 7026 39136 7042 39200
rect 7106 39136 7122 39200
rect 7186 39136 7194 39200
rect 6874 39135 7194 39136
rect 12805 39200 13125 39201
rect 12805 39136 12813 39200
rect 12877 39136 12893 39200
rect 12957 39136 12973 39200
rect 13037 39136 13053 39200
rect 13117 39136 13125 39200
rect 12805 39135 13125 39136
rect 3909 38656 4229 38657
rect 3909 38592 3917 38656
rect 3981 38592 3997 38656
rect 4061 38592 4077 38656
rect 4141 38592 4157 38656
rect 4221 38592 4229 38656
rect 3909 38591 4229 38592
rect 9840 38656 10160 38657
rect 9840 38592 9848 38656
rect 9912 38592 9928 38656
rect 9992 38592 10008 38656
rect 10072 38592 10088 38656
rect 10152 38592 10160 38656
rect 9840 38591 10160 38592
rect 15770 38656 16090 38657
rect 15770 38592 15778 38656
rect 15842 38592 15858 38656
rect 15922 38592 15938 38656
rect 16002 38592 16018 38656
rect 16082 38592 16090 38656
rect 15770 38591 16090 38592
rect 6874 38112 7194 38113
rect 6874 38048 6882 38112
rect 6946 38048 6962 38112
rect 7026 38048 7042 38112
rect 7106 38048 7122 38112
rect 7186 38048 7194 38112
rect 6874 38047 7194 38048
rect 12805 38112 13125 38113
rect 12805 38048 12813 38112
rect 12877 38048 12893 38112
rect 12957 38048 12973 38112
rect 13037 38048 13053 38112
rect 13117 38048 13125 38112
rect 12805 38047 13125 38048
rect 3909 37568 4229 37569
rect 3909 37504 3917 37568
rect 3981 37504 3997 37568
rect 4061 37504 4077 37568
rect 4141 37504 4157 37568
rect 4221 37504 4229 37568
rect 3909 37503 4229 37504
rect 9840 37568 10160 37569
rect 9840 37504 9848 37568
rect 9912 37504 9928 37568
rect 9992 37504 10008 37568
rect 10072 37504 10088 37568
rect 10152 37504 10160 37568
rect 9840 37503 10160 37504
rect 15770 37568 16090 37569
rect 15770 37504 15778 37568
rect 15842 37504 15858 37568
rect 15922 37504 15938 37568
rect 16002 37504 16018 37568
rect 16082 37504 16090 37568
rect 15770 37503 16090 37504
rect 6874 37024 7194 37025
rect 6874 36960 6882 37024
rect 6946 36960 6962 37024
rect 7026 36960 7042 37024
rect 7106 36960 7122 37024
rect 7186 36960 7194 37024
rect 6874 36959 7194 36960
rect 12805 37024 13125 37025
rect 12805 36960 12813 37024
rect 12877 36960 12893 37024
rect 12957 36960 12973 37024
rect 13037 36960 13053 37024
rect 13117 36960 13125 37024
rect 12805 36959 13125 36960
rect 3909 36480 4229 36481
rect 3909 36416 3917 36480
rect 3981 36416 3997 36480
rect 4061 36416 4077 36480
rect 4141 36416 4157 36480
rect 4221 36416 4229 36480
rect 3909 36415 4229 36416
rect 9840 36480 10160 36481
rect 9840 36416 9848 36480
rect 9912 36416 9928 36480
rect 9992 36416 10008 36480
rect 10072 36416 10088 36480
rect 10152 36416 10160 36480
rect 9840 36415 10160 36416
rect 15770 36480 16090 36481
rect 15770 36416 15778 36480
rect 15842 36416 15858 36480
rect 15922 36416 15938 36480
rect 16002 36416 16018 36480
rect 16082 36416 16090 36480
rect 15770 36415 16090 36416
rect 0 36138 800 36168
rect 1853 36138 1919 36141
rect 0 36136 1919 36138
rect 0 36080 1858 36136
rect 1914 36080 1919 36136
rect 0 36078 1919 36080
rect 0 36048 800 36078
rect 1853 36075 1919 36078
rect 6874 35936 7194 35937
rect 6874 35872 6882 35936
rect 6946 35872 6962 35936
rect 7026 35872 7042 35936
rect 7106 35872 7122 35936
rect 7186 35872 7194 35936
rect 6874 35871 7194 35872
rect 12805 35936 13125 35937
rect 12805 35872 12813 35936
rect 12877 35872 12893 35936
rect 12957 35872 12973 35936
rect 13037 35872 13053 35936
rect 13117 35872 13125 35936
rect 12805 35871 13125 35872
rect 3909 35392 4229 35393
rect 3909 35328 3917 35392
rect 3981 35328 3997 35392
rect 4061 35328 4077 35392
rect 4141 35328 4157 35392
rect 4221 35328 4229 35392
rect 3909 35327 4229 35328
rect 9840 35392 10160 35393
rect 9840 35328 9848 35392
rect 9912 35328 9928 35392
rect 9992 35328 10008 35392
rect 10072 35328 10088 35392
rect 10152 35328 10160 35392
rect 9840 35327 10160 35328
rect 15770 35392 16090 35393
rect 15770 35328 15778 35392
rect 15842 35328 15858 35392
rect 15922 35328 15938 35392
rect 16002 35328 16018 35392
rect 16082 35328 16090 35392
rect 15770 35327 16090 35328
rect 6874 34848 7194 34849
rect 6874 34784 6882 34848
rect 6946 34784 6962 34848
rect 7026 34784 7042 34848
rect 7106 34784 7122 34848
rect 7186 34784 7194 34848
rect 6874 34783 7194 34784
rect 12805 34848 13125 34849
rect 12805 34784 12813 34848
rect 12877 34784 12893 34848
rect 12957 34784 12973 34848
rect 13037 34784 13053 34848
rect 13117 34784 13125 34848
rect 12805 34783 13125 34784
rect 15745 34642 15811 34645
rect 16941 34642 17007 34645
rect 15745 34640 17007 34642
rect 15745 34584 15750 34640
rect 15806 34584 16946 34640
rect 17002 34584 17007 34640
rect 15745 34582 17007 34584
rect 15745 34579 15811 34582
rect 16941 34579 17007 34582
rect 15653 34506 15719 34509
rect 19200 34506 20000 34536
rect 15653 34504 20000 34506
rect 15653 34448 15658 34504
rect 15714 34448 20000 34504
rect 15653 34446 20000 34448
rect 15653 34443 15719 34446
rect 19200 34416 20000 34446
rect 3909 34304 4229 34305
rect 3909 34240 3917 34304
rect 3981 34240 3997 34304
rect 4061 34240 4077 34304
rect 4141 34240 4157 34304
rect 4221 34240 4229 34304
rect 3909 34239 4229 34240
rect 9840 34304 10160 34305
rect 9840 34240 9848 34304
rect 9912 34240 9928 34304
rect 9992 34240 10008 34304
rect 10072 34240 10088 34304
rect 10152 34240 10160 34304
rect 9840 34239 10160 34240
rect 15770 34304 16090 34305
rect 15770 34240 15778 34304
rect 15842 34240 15858 34304
rect 15922 34240 15938 34304
rect 16002 34240 16018 34304
rect 16082 34240 16090 34304
rect 15770 34239 16090 34240
rect 6874 33760 7194 33761
rect 6874 33696 6882 33760
rect 6946 33696 6962 33760
rect 7026 33696 7042 33760
rect 7106 33696 7122 33760
rect 7186 33696 7194 33760
rect 6874 33695 7194 33696
rect 12805 33760 13125 33761
rect 12805 33696 12813 33760
rect 12877 33696 12893 33760
rect 12957 33696 12973 33760
rect 13037 33696 13053 33760
rect 13117 33696 13125 33760
rect 12805 33695 13125 33696
rect 13537 33554 13603 33557
rect 15561 33554 15627 33557
rect 17585 33554 17651 33557
rect 13537 33552 17651 33554
rect 13537 33496 13542 33552
rect 13598 33496 15566 33552
rect 15622 33496 17590 33552
rect 17646 33496 17651 33552
rect 13537 33494 17651 33496
rect 13537 33491 13603 33494
rect 15561 33491 15627 33494
rect 17585 33491 17651 33494
rect 16573 33284 16639 33285
rect 16573 33280 16620 33284
rect 16684 33282 16690 33284
rect 16573 33224 16578 33280
rect 16573 33220 16620 33224
rect 16684 33222 16730 33282
rect 16684 33220 16690 33222
rect 16573 33219 16639 33220
rect 3909 33216 4229 33217
rect 3909 33152 3917 33216
rect 3981 33152 3997 33216
rect 4061 33152 4077 33216
rect 4141 33152 4157 33216
rect 4221 33152 4229 33216
rect 3909 33151 4229 33152
rect 9840 33216 10160 33217
rect 9840 33152 9848 33216
rect 9912 33152 9928 33216
rect 9992 33152 10008 33216
rect 10072 33152 10088 33216
rect 10152 33152 10160 33216
rect 9840 33151 10160 33152
rect 15770 33216 16090 33217
rect 15770 33152 15778 33216
rect 15842 33152 15858 33216
rect 15922 33152 15938 33216
rect 16002 33152 16018 33216
rect 16082 33152 16090 33216
rect 15770 33151 16090 33152
rect 6874 32672 7194 32673
rect 6874 32608 6882 32672
rect 6946 32608 6962 32672
rect 7026 32608 7042 32672
rect 7106 32608 7122 32672
rect 7186 32608 7194 32672
rect 6874 32607 7194 32608
rect 12805 32672 13125 32673
rect 12805 32608 12813 32672
rect 12877 32608 12893 32672
rect 12957 32608 12973 32672
rect 13037 32608 13053 32672
rect 13117 32608 13125 32672
rect 12805 32607 13125 32608
rect 3909 32128 4229 32129
rect 3909 32064 3917 32128
rect 3981 32064 3997 32128
rect 4061 32064 4077 32128
rect 4141 32064 4157 32128
rect 4221 32064 4229 32128
rect 3909 32063 4229 32064
rect 9840 32128 10160 32129
rect 9840 32064 9848 32128
rect 9912 32064 9928 32128
rect 9992 32064 10008 32128
rect 10072 32064 10088 32128
rect 10152 32064 10160 32128
rect 9840 32063 10160 32064
rect 15770 32128 16090 32129
rect 15770 32064 15778 32128
rect 15842 32064 15858 32128
rect 15922 32064 15938 32128
rect 16002 32064 16018 32128
rect 16082 32064 16090 32128
rect 15770 32063 16090 32064
rect 6874 31584 7194 31585
rect 6874 31520 6882 31584
rect 6946 31520 6962 31584
rect 7026 31520 7042 31584
rect 7106 31520 7122 31584
rect 7186 31520 7194 31584
rect 6874 31519 7194 31520
rect 12805 31584 13125 31585
rect 12805 31520 12813 31584
rect 12877 31520 12893 31584
rect 12957 31520 12973 31584
rect 13037 31520 13053 31584
rect 13117 31520 13125 31584
rect 12805 31519 13125 31520
rect 3909 31040 4229 31041
rect 3909 30976 3917 31040
rect 3981 30976 3997 31040
rect 4061 30976 4077 31040
rect 4141 30976 4157 31040
rect 4221 30976 4229 31040
rect 3909 30975 4229 30976
rect 9840 31040 10160 31041
rect 9840 30976 9848 31040
rect 9912 30976 9928 31040
rect 9992 30976 10008 31040
rect 10072 30976 10088 31040
rect 10152 30976 10160 31040
rect 9840 30975 10160 30976
rect 15770 31040 16090 31041
rect 15770 30976 15778 31040
rect 15842 30976 15858 31040
rect 15922 30976 15938 31040
rect 16002 30976 16018 31040
rect 16082 30976 16090 31040
rect 15770 30975 16090 30976
rect 0 30562 800 30592
rect 1393 30562 1459 30565
rect 0 30560 1459 30562
rect 0 30504 1398 30560
rect 1454 30504 1459 30560
rect 0 30502 1459 30504
rect 0 30472 800 30502
rect 1393 30499 1459 30502
rect 6874 30496 7194 30497
rect 6874 30432 6882 30496
rect 6946 30432 6962 30496
rect 7026 30432 7042 30496
rect 7106 30432 7122 30496
rect 7186 30432 7194 30496
rect 6874 30431 7194 30432
rect 12805 30496 13125 30497
rect 12805 30432 12813 30496
rect 12877 30432 12893 30496
rect 12957 30432 12973 30496
rect 13037 30432 13053 30496
rect 13117 30432 13125 30496
rect 12805 30431 13125 30432
rect 3909 29952 4229 29953
rect 3909 29888 3917 29952
rect 3981 29888 3997 29952
rect 4061 29888 4077 29952
rect 4141 29888 4157 29952
rect 4221 29888 4229 29952
rect 3909 29887 4229 29888
rect 9840 29952 10160 29953
rect 9840 29888 9848 29952
rect 9912 29888 9928 29952
rect 9992 29888 10008 29952
rect 10072 29888 10088 29952
rect 10152 29888 10160 29952
rect 9840 29887 10160 29888
rect 15770 29952 16090 29953
rect 15770 29888 15778 29952
rect 15842 29888 15858 29952
rect 15922 29888 15938 29952
rect 16002 29888 16018 29952
rect 16082 29888 16090 29952
rect 15770 29887 16090 29888
rect 6874 29408 7194 29409
rect 6874 29344 6882 29408
rect 6946 29344 6962 29408
rect 7026 29344 7042 29408
rect 7106 29344 7122 29408
rect 7186 29344 7194 29408
rect 6874 29343 7194 29344
rect 12805 29408 13125 29409
rect 12805 29344 12813 29408
rect 12877 29344 12893 29408
rect 12957 29344 12973 29408
rect 13037 29344 13053 29408
rect 13117 29344 13125 29408
rect 12805 29343 13125 29344
rect 3909 28864 4229 28865
rect 3909 28800 3917 28864
rect 3981 28800 3997 28864
rect 4061 28800 4077 28864
rect 4141 28800 4157 28864
rect 4221 28800 4229 28864
rect 3909 28799 4229 28800
rect 9840 28864 10160 28865
rect 9840 28800 9848 28864
rect 9912 28800 9928 28864
rect 9992 28800 10008 28864
rect 10072 28800 10088 28864
rect 10152 28800 10160 28864
rect 9840 28799 10160 28800
rect 15770 28864 16090 28865
rect 15770 28800 15778 28864
rect 15842 28800 15858 28864
rect 15922 28800 15938 28864
rect 16002 28800 16018 28864
rect 16082 28800 16090 28864
rect 15770 28799 16090 28800
rect 6874 28320 7194 28321
rect 6874 28256 6882 28320
rect 6946 28256 6962 28320
rect 7026 28256 7042 28320
rect 7106 28256 7122 28320
rect 7186 28256 7194 28320
rect 6874 28255 7194 28256
rect 12805 28320 13125 28321
rect 12805 28256 12813 28320
rect 12877 28256 12893 28320
rect 12957 28256 12973 28320
rect 13037 28256 13053 28320
rect 13117 28256 13125 28320
rect 12805 28255 13125 28256
rect 18137 28250 18203 28253
rect 19200 28250 20000 28280
rect 18137 28248 20000 28250
rect 18137 28192 18142 28248
rect 18198 28192 20000 28248
rect 18137 28190 20000 28192
rect 18137 28187 18203 28190
rect 19200 28160 20000 28190
rect 3909 27776 4229 27777
rect 3909 27712 3917 27776
rect 3981 27712 3997 27776
rect 4061 27712 4077 27776
rect 4141 27712 4157 27776
rect 4221 27712 4229 27776
rect 3909 27711 4229 27712
rect 9840 27776 10160 27777
rect 9840 27712 9848 27776
rect 9912 27712 9928 27776
rect 9992 27712 10008 27776
rect 10072 27712 10088 27776
rect 10152 27712 10160 27776
rect 9840 27711 10160 27712
rect 15770 27776 16090 27777
rect 15770 27712 15778 27776
rect 15842 27712 15858 27776
rect 15922 27712 15938 27776
rect 16002 27712 16018 27776
rect 16082 27712 16090 27776
rect 15770 27711 16090 27712
rect 6874 27232 7194 27233
rect 6874 27168 6882 27232
rect 6946 27168 6962 27232
rect 7026 27168 7042 27232
rect 7106 27168 7122 27232
rect 7186 27168 7194 27232
rect 6874 27167 7194 27168
rect 12805 27232 13125 27233
rect 12805 27168 12813 27232
rect 12877 27168 12893 27232
rect 12957 27168 12973 27232
rect 13037 27168 13053 27232
rect 13117 27168 13125 27232
rect 12805 27167 13125 27168
rect 3909 26688 4229 26689
rect 3909 26624 3917 26688
rect 3981 26624 3997 26688
rect 4061 26624 4077 26688
rect 4141 26624 4157 26688
rect 4221 26624 4229 26688
rect 3909 26623 4229 26624
rect 9840 26688 10160 26689
rect 9840 26624 9848 26688
rect 9912 26624 9928 26688
rect 9992 26624 10008 26688
rect 10072 26624 10088 26688
rect 10152 26624 10160 26688
rect 9840 26623 10160 26624
rect 15770 26688 16090 26689
rect 15770 26624 15778 26688
rect 15842 26624 15858 26688
rect 15922 26624 15938 26688
rect 16002 26624 16018 26688
rect 16082 26624 16090 26688
rect 15770 26623 16090 26624
rect 6874 26144 7194 26145
rect 6874 26080 6882 26144
rect 6946 26080 6962 26144
rect 7026 26080 7042 26144
rect 7106 26080 7122 26144
rect 7186 26080 7194 26144
rect 6874 26079 7194 26080
rect 12805 26144 13125 26145
rect 12805 26080 12813 26144
rect 12877 26080 12893 26144
rect 12957 26080 12973 26144
rect 13037 26080 13053 26144
rect 13117 26080 13125 26144
rect 12805 26079 13125 26080
rect 3909 25600 4229 25601
rect 3909 25536 3917 25600
rect 3981 25536 3997 25600
rect 4061 25536 4077 25600
rect 4141 25536 4157 25600
rect 4221 25536 4229 25600
rect 3909 25535 4229 25536
rect 9840 25600 10160 25601
rect 9840 25536 9848 25600
rect 9912 25536 9928 25600
rect 9992 25536 10008 25600
rect 10072 25536 10088 25600
rect 10152 25536 10160 25600
rect 9840 25535 10160 25536
rect 15770 25600 16090 25601
rect 15770 25536 15778 25600
rect 15842 25536 15858 25600
rect 15922 25536 15938 25600
rect 16002 25536 16018 25600
rect 16082 25536 16090 25600
rect 15770 25535 16090 25536
rect 13169 25530 13235 25533
rect 15510 25530 15516 25532
rect 13169 25528 15516 25530
rect 13169 25472 13174 25528
rect 13230 25472 15516 25528
rect 13169 25470 15516 25472
rect 13169 25467 13235 25470
rect 15510 25468 15516 25470
rect 15580 25468 15586 25532
rect 6874 25056 7194 25057
rect 0 24986 800 25016
rect 6874 24992 6882 25056
rect 6946 24992 6962 25056
rect 7026 24992 7042 25056
rect 7106 24992 7122 25056
rect 7186 24992 7194 25056
rect 6874 24991 7194 24992
rect 12805 25056 13125 25057
rect 12805 24992 12813 25056
rect 12877 24992 12893 25056
rect 12957 24992 12973 25056
rect 13037 24992 13053 25056
rect 13117 24992 13125 25056
rect 12805 24991 13125 24992
rect 1485 24986 1551 24989
rect 0 24984 1551 24986
rect 0 24928 1490 24984
rect 1546 24928 1551 24984
rect 0 24926 1551 24928
rect 0 24896 800 24926
rect 1485 24923 1551 24926
rect 3909 24512 4229 24513
rect 3909 24448 3917 24512
rect 3981 24448 3997 24512
rect 4061 24448 4077 24512
rect 4141 24448 4157 24512
rect 4221 24448 4229 24512
rect 3909 24447 4229 24448
rect 9840 24512 10160 24513
rect 9840 24448 9848 24512
rect 9912 24448 9928 24512
rect 9992 24448 10008 24512
rect 10072 24448 10088 24512
rect 10152 24448 10160 24512
rect 9840 24447 10160 24448
rect 15770 24512 16090 24513
rect 15770 24448 15778 24512
rect 15842 24448 15858 24512
rect 15922 24448 15938 24512
rect 16002 24448 16018 24512
rect 16082 24448 16090 24512
rect 15770 24447 16090 24448
rect 6874 23968 7194 23969
rect 6874 23904 6882 23968
rect 6946 23904 6962 23968
rect 7026 23904 7042 23968
rect 7106 23904 7122 23968
rect 7186 23904 7194 23968
rect 6874 23903 7194 23904
rect 12805 23968 13125 23969
rect 12805 23904 12813 23968
rect 12877 23904 12893 23968
rect 12957 23904 12973 23968
rect 13037 23904 13053 23968
rect 13117 23904 13125 23968
rect 12805 23903 13125 23904
rect 3909 23424 4229 23425
rect 3909 23360 3917 23424
rect 3981 23360 3997 23424
rect 4061 23360 4077 23424
rect 4141 23360 4157 23424
rect 4221 23360 4229 23424
rect 3909 23359 4229 23360
rect 9840 23424 10160 23425
rect 9840 23360 9848 23424
rect 9912 23360 9928 23424
rect 9992 23360 10008 23424
rect 10072 23360 10088 23424
rect 10152 23360 10160 23424
rect 9840 23359 10160 23360
rect 15770 23424 16090 23425
rect 15770 23360 15778 23424
rect 15842 23360 15858 23424
rect 15922 23360 15938 23424
rect 16002 23360 16018 23424
rect 16082 23360 16090 23424
rect 15770 23359 16090 23360
rect 6874 22880 7194 22881
rect 6874 22816 6882 22880
rect 6946 22816 6962 22880
rect 7026 22816 7042 22880
rect 7106 22816 7122 22880
rect 7186 22816 7194 22880
rect 6874 22815 7194 22816
rect 12805 22880 13125 22881
rect 12805 22816 12813 22880
rect 12877 22816 12893 22880
rect 12957 22816 12973 22880
rect 13037 22816 13053 22880
rect 13117 22816 13125 22880
rect 12805 22815 13125 22816
rect 3909 22336 4229 22337
rect 3909 22272 3917 22336
rect 3981 22272 3997 22336
rect 4061 22272 4077 22336
rect 4141 22272 4157 22336
rect 4221 22272 4229 22336
rect 3909 22271 4229 22272
rect 9840 22336 10160 22337
rect 9840 22272 9848 22336
rect 9912 22272 9928 22336
rect 9992 22272 10008 22336
rect 10072 22272 10088 22336
rect 10152 22272 10160 22336
rect 9840 22271 10160 22272
rect 15770 22336 16090 22337
rect 15770 22272 15778 22336
rect 15842 22272 15858 22336
rect 15922 22272 15938 22336
rect 16002 22272 16018 22336
rect 16082 22272 16090 22336
rect 15770 22271 16090 22272
rect 18137 21994 18203 21997
rect 19200 21994 20000 22024
rect 18137 21992 20000 21994
rect 18137 21936 18142 21992
rect 18198 21936 20000 21992
rect 18137 21934 20000 21936
rect 18137 21931 18203 21934
rect 19200 21904 20000 21934
rect 6874 21792 7194 21793
rect 6874 21728 6882 21792
rect 6946 21728 6962 21792
rect 7026 21728 7042 21792
rect 7106 21728 7122 21792
rect 7186 21728 7194 21792
rect 6874 21727 7194 21728
rect 12805 21792 13125 21793
rect 12805 21728 12813 21792
rect 12877 21728 12893 21792
rect 12957 21728 12973 21792
rect 13037 21728 13053 21792
rect 13117 21728 13125 21792
rect 12805 21727 13125 21728
rect 3909 21248 4229 21249
rect 3909 21184 3917 21248
rect 3981 21184 3997 21248
rect 4061 21184 4077 21248
rect 4141 21184 4157 21248
rect 4221 21184 4229 21248
rect 3909 21183 4229 21184
rect 9840 21248 10160 21249
rect 9840 21184 9848 21248
rect 9912 21184 9928 21248
rect 9992 21184 10008 21248
rect 10072 21184 10088 21248
rect 10152 21184 10160 21248
rect 9840 21183 10160 21184
rect 15770 21248 16090 21249
rect 15770 21184 15778 21248
rect 15842 21184 15858 21248
rect 15922 21184 15938 21248
rect 16002 21184 16018 21248
rect 16082 21184 16090 21248
rect 15770 21183 16090 21184
rect 6874 20704 7194 20705
rect 6874 20640 6882 20704
rect 6946 20640 6962 20704
rect 7026 20640 7042 20704
rect 7106 20640 7122 20704
rect 7186 20640 7194 20704
rect 6874 20639 7194 20640
rect 12805 20704 13125 20705
rect 12805 20640 12813 20704
rect 12877 20640 12893 20704
rect 12957 20640 12973 20704
rect 13037 20640 13053 20704
rect 13117 20640 13125 20704
rect 12805 20639 13125 20640
rect 3909 20160 4229 20161
rect 3909 20096 3917 20160
rect 3981 20096 3997 20160
rect 4061 20096 4077 20160
rect 4141 20096 4157 20160
rect 4221 20096 4229 20160
rect 3909 20095 4229 20096
rect 9840 20160 10160 20161
rect 9840 20096 9848 20160
rect 9912 20096 9928 20160
rect 9992 20096 10008 20160
rect 10072 20096 10088 20160
rect 10152 20096 10160 20160
rect 9840 20095 10160 20096
rect 15770 20160 16090 20161
rect 15770 20096 15778 20160
rect 15842 20096 15858 20160
rect 15922 20096 15938 20160
rect 16002 20096 16018 20160
rect 16082 20096 16090 20160
rect 15770 20095 16090 20096
rect 6874 19616 7194 19617
rect 6874 19552 6882 19616
rect 6946 19552 6962 19616
rect 7026 19552 7042 19616
rect 7106 19552 7122 19616
rect 7186 19552 7194 19616
rect 6874 19551 7194 19552
rect 12805 19616 13125 19617
rect 12805 19552 12813 19616
rect 12877 19552 12893 19616
rect 12957 19552 12973 19616
rect 13037 19552 13053 19616
rect 13117 19552 13125 19616
rect 12805 19551 13125 19552
rect 0 19410 800 19440
rect 1393 19410 1459 19413
rect 0 19408 1459 19410
rect 0 19352 1398 19408
rect 1454 19352 1459 19408
rect 0 19350 1459 19352
rect 0 19320 800 19350
rect 1393 19347 1459 19350
rect 3909 19072 4229 19073
rect 3909 19008 3917 19072
rect 3981 19008 3997 19072
rect 4061 19008 4077 19072
rect 4141 19008 4157 19072
rect 4221 19008 4229 19072
rect 3909 19007 4229 19008
rect 9840 19072 10160 19073
rect 9840 19008 9848 19072
rect 9912 19008 9928 19072
rect 9992 19008 10008 19072
rect 10072 19008 10088 19072
rect 10152 19008 10160 19072
rect 9840 19007 10160 19008
rect 15770 19072 16090 19073
rect 15770 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15938 19072
rect 16002 19008 16018 19072
rect 16082 19008 16090 19072
rect 15770 19007 16090 19008
rect 6874 18528 7194 18529
rect 6874 18464 6882 18528
rect 6946 18464 6962 18528
rect 7026 18464 7042 18528
rect 7106 18464 7122 18528
rect 7186 18464 7194 18528
rect 6874 18463 7194 18464
rect 12805 18528 13125 18529
rect 12805 18464 12813 18528
rect 12877 18464 12893 18528
rect 12957 18464 12973 18528
rect 13037 18464 13053 18528
rect 13117 18464 13125 18528
rect 12805 18463 13125 18464
rect 3909 17984 4229 17985
rect 3909 17920 3917 17984
rect 3981 17920 3997 17984
rect 4061 17920 4077 17984
rect 4141 17920 4157 17984
rect 4221 17920 4229 17984
rect 3909 17919 4229 17920
rect 9840 17984 10160 17985
rect 9840 17920 9848 17984
rect 9912 17920 9928 17984
rect 9992 17920 10008 17984
rect 10072 17920 10088 17984
rect 10152 17920 10160 17984
rect 9840 17919 10160 17920
rect 15770 17984 16090 17985
rect 15770 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15938 17984
rect 16002 17920 16018 17984
rect 16082 17920 16090 17984
rect 15770 17919 16090 17920
rect 6874 17440 7194 17441
rect 6874 17376 6882 17440
rect 6946 17376 6962 17440
rect 7026 17376 7042 17440
rect 7106 17376 7122 17440
rect 7186 17376 7194 17440
rect 6874 17375 7194 17376
rect 12805 17440 13125 17441
rect 12805 17376 12813 17440
rect 12877 17376 12893 17440
rect 12957 17376 12973 17440
rect 13037 17376 13053 17440
rect 13117 17376 13125 17440
rect 12805 17375 13125 17376
rect 3909 16896 4229 16897
rect 3909 16832 3917 16896
rect 3981 16832 3997 16896
rect 4061 16832 4077 16896
rect 4141 16832 4157 16896
rect 4221 16832 4229 16896
rect 3909 16831 4229 16832
rect 9840 16896 10160 16897
rect 9840 16832 9848 16896
rect 9912 16832 9928 16896
rect 9992 16832 10008 16896
rect 10072 16832 10088 16896
rect 10152 16832 10160 16896
rect 9840 16831 10160 16832
rect 15770 16896 16090 16897
rect 15770 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15938 16896
rect 16002 16832 16018 16896
rect 16082 16832 16090 16896
rect 15770 16831 16090 16832
rect 6874 16352 7194 16353
rect 6874 16288 6882 16352
rect 6946 16288 6962 16352
rect 7026 16288 7042 16352
rect 7106 16288 7122 16352
rect 7186 16288 7194 16352
rect 6874 16287 7194 16288
rect 12805 16352 13125 16353
rect 12805 16288 12813 16352
rect 12877 16288 12893 16352
rect 12957 16288 12973 16352
rect 13037 16288 13053 16352
rect 13117 16288 13125 16352
rect 12805 16287 13125 16288
rect 3909 15808 4229 15809
rect 3909 15744 3917 15808
rect 3981 15744 3997 15808
rect 4061 15744 4077 15808
rect 4141 15744 4157 15808
rect 4221 15744 4229 15808
rect 3909 15743 4229 15744
rect 9840 15808 10160 15809
rect 9840 15744 9848 15808
rect 9912 15744 9928 15808
rect 9992 15744 10008 15808
rect 10072 15744 10088 15808
rect 10152 15744 10160 15808
rect 9840 15743 10160 15744
rect 15770 15808 16090 15809
rect 15770 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15938 15808
rect 16002 15744 16018 15808
rect 16082 15744 16090 15808
rect 15770 15743 16090 15744
rect 18137 15738 18203 15741
rect 19200 15738 20000 15768
rect 18137 15736 20000 15738
rect 18137 15680 18142 15736
rect 18198 15680 20000 15736
rect 18137 15678 20000 15680
rect 18137 15675 18203 15678
rect 19200 15648 20000 15678
rect 6874 15264 7194 15265
rect 6874 15200 6882 15264
rect 6946 15200 6962 15264
rect 7026 15200 7042 15264
rect 7106 15200 7122 15264
rect 7186 15200 7194 15264
rect 6874 15199 7194 15200
rect 12805 15264 13125 15265
rect 12805 15200 12813 15264
rect 12877 15200 12893 15264
rect 12957 15200 12973 15264
rect 13037 15200 13053 15264
rect 13117 15200 13125 15264
rect 12805 15199 13125 15200
rect 3909 14720 4229 14721
rect 3909 14656 3917 14720
rect 3981 14656 3997 14720
rect 4061 14656 4077 14720
rect 4141 14656 4157 14720
rect 4221 14656 4229 14720
rect 3909 14655 4229 14656
rect 9840 14720 10160 14721
rect 9840 14656 9848 14720
rect 9912 14656 9928 14720
rect 9992 14656 10008 14720
rect 10072 14656 10088 14720
rect 10152 14656 10160 14720
rect 9840 14655 10160 14656
rect 15770 14720 16090 14721
rect 15770 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15938 14720
rect 16002 14656 16018 14720
rect 16082 14656 16090 14720
rect 15770 14655 16090 14656
rect 6874 14176 7194 14177
rect 6874 14112 6882 14176
rect 6946 14112 6962 14176
rect 7026 14112 7042 14176
rect 7106 14112 7122 14176
rect 7186 14112 7194 14176
rect 6874 14111 7194 14112
rect 12805 14176 13125 14177
rect 12805 14112 12813 14176
rect 12877 14112 12893 14176
rect 12957 14112 12973 14176
rect 13037 14112 13053 14176
rect 13117 14112 13125 14176
rect 12805 14111 13125 14112
rect 0 13834 800 13864
rect 1393 13834 1459 13837
rect 0 13832 1459 13834
rect 0 13776 1398 13832
rect 1454 13776 1459 13832
rect 0 13774 1459 13776
rect 0 13744 800 13774
rect 1393 13771 1459 13774
rect 3909 13632 4229 13633
rect 3909 13568 3917 13632
rect 3981 13568 3997 13632
rect 4061 13568 4077 13632
rect 4141 13568 4157 13632
rect 4221 13568 4229 13632
rect 3909 13567 4229 13568
rect 9840 13632 10160 13633
rect 9840 13568 9848 13632
rect 9912 13568 9928 13632
rect 9992 13568 10008 13632
rect 10072 13568 10088 13632
rect 10152 13568 10160 13632
rect 9840 13567 10160 13568
rect 15770 13632 16090 13633
rect 15770 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15938 13632
rect 16002 13568 16018 13632
rect 16082 13568 16090 13632
rect 15770 13567 16090 13568
rect 6874 13088 7194 13089
rect 6874 13024 6882 13088
rect 6946 13024 6962 13088
rect 7026 13024 7042 13088
rect 7106 13024 7122 13088
rect 7186 13024 7194 13088
rect 6874 13023 7194 13024
rect 12805 13088 13125 13089
rect 12805 13024 12813 13088
rect 12877 13024 12893 13088
rect 12957 13024 12973 13088
rect 13037 13024 13053 13088
rect 13117 13024 13125 13088
rect 12805 13023 13125 13024
rect 3909 12544 4229 12545
rect 3909 12480 3917 12544
rect 3981 12480 3997 12544
rect 4061 12480 4077 12544
rect 4141 12480 4157 12544
rect 4221 12480 4229 12544
rect 3909 12479 4229 12480
rect 9840 12544 10160 12545
rect 9840 12480 9848 12544
rect 9912 12480 9928 12544
rect 9992 12480 10008 12544
rect 10072 12480 10088 12544
rect 10152 12480 10160 12544
rect 9840 12479 10160 12480
rect 15770 12544 16090 12545
rect 15770 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15938 12544
rect 16002 12480 16018 12544
rect 16082 12480 16090 12544
rect 15770 12479 16090 12480
rect 6874 12000 7194 12001
rect 6874 11936 6882 12000
rect 6946 11936 6962 12000
rect 7026 11936 7042 12000
rect 7106 11936 7122 12000
rect 7186 11936 7194 12000
rect 6874 11935 7194 11936
rect 12805 12000 13125 12001
rect 12805 11936 12813 12000
rect 12877 11936 12893 12000
rect 12957 11936 12973 12000
rect 13037 11936 13053 12000
rect 13117 11936 13125 12000
rect 12805 11935 13125 11936
rect 3909 11456 4229 11457
rect 3909 11392 3917 11456
rect 3981 11392 3997 11456
rect 4061 11392 4077 11456
rect 4141 11392 4157 11456
rect 4221 11392 4229 11456
rect 3909 11391 4229 11392
rect 9840 11456 10160 11457
rect 9840 11392 9848 11456
rect 9912 11392 9928 11456
rect 9992 11392 10008 11456
rect 10072 11392 10088 11456
rect 10152 11392 10160 11456
rect 9840 11391 10160 11392
rect 15770 11456 16090 11457
rect 15770 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15938 11456
rect 16002 11392 16018 11456
rect 16082 11392 16090 11456
rect 15770 11391 16090 11392
rect 6874 10912 7194 10913
rect 6874 10848 6882 10912
rect 6946 10848 6962 10912
rect 7026 10848 7042 10912
rect 7106 10848 7122 10912
rect 7186 10848 7194 10912
rect 6874 10847 7194 10848
rect 12805 10912 13125 10913
rect 12805 10848 12813 10912
rect 12877 10848 12893 10912
rect 12957 10848 12973 10912
rect 13037 10848 13053 10912
rect 13117 10848 13125 10912
rect 12805 10847 13125 10848
rect 3909 10368 4229 10369
rect 3909 10304 3917 10368
rect 3981 10304 3997 10368
rect 4061 10304 4077 10368
rect 4141 10304 4157 10368
rect 4221 10304 4229 10368
rect 3909 10303 4229 10304
rect 9840 10368 10160 10369
rect 9840 10304 9848 10368
rect 9912 10304 9928 10368
rect 9992 10304 10008 10368
rect 10072 10304 10088 10368
rect 10152 10304 10160 10368
rect 9840 10303 10160 10304
rect 15770 10368 16090 10369
rect 15770 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15938 10368
rect 16002 10304 16018 10368
rect 16082 10304 16090 10368
rect 15770 10303 16090 10304
rect 6874 9824 7194 9825
rect 6874 9760 6882 9824
rect 6946 9760 6962 9824
rect 7026 9760 7042 9824
rect 7106 9760 7122 9824
rect 7186 9760 7194 9824
rect 6874 9759 7194 9760
rect 12805 9824 13125 9825
rect 12805 9760 12813 9824
rect 12877 9760 12893 9824
rect 12957 9760 12973 9824
rect 13037 9760 13053 9824
rect 13117 9760 13125 9824
rect 12805 9759 13125 9760
rect 18045 9482 18111 9485
rect 19200 9482 20000 9512
rect 18045 9480 20000 9482
rect 18045 9424 18050 9480
rect 18106 9424 20000 9480
rect 18045 9422 20000 9424
rect 18045 9419 18111 9422
rect 19200 9392 20000 9422
rect 3909 9280 4229 9281
rect 3909 9216 3917 9280
rect 3981 9216 3997 9280
rect 4061 9216 4077 9280
rect 4141 9216 4157 9280
rect 4221 9216 4229 9280
rect 3909 9215 4229 9216
rect 9840 9280 10160 9281
rect 9840 9216 9848 9280
rect 9912 9216 9928 9280
rect 9992 9216 10008 9280
rect 10072 9216 10088 9280
rect 10152 9216 10160 9280
rect 9840 9215 10160 9216
rect 15770 9280 16090 9281
rect 15770 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15938 9280
rect 16002 9216 16018 9280
rect 16082 9216 16090 9280
rect 15770 9215 16090 9216
rect 6874 8736 7194 8737
rect 6874 8672 6882 8736
rect 6946 8672 6962 8736
rect 7026 8672 7042 8736
rect 7106 8672 7122 8736
rect 7186 8672 7194 8736
rect 6874 8671 7194 8672
rect 12805 8736 13125 8737
rect 12805 8672 12813 8736
rect 12877 8672 12893 8736
rect 12957 8672 12973 8736
rect 13037 8672 13053 8736
rect 13117 8672 13125 8736
rect 12805 8671 13125 8672
rect 0 8258 800 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 800 8198
rect 1577 8195 1643 8198
rect 3909 8192 4229 8193
rect 3909 8128 3917 8192
rect 3981 8128 3997 8192
rect 4061 8128 4077 8192
rect 4141 8128 4157 8192
rect 4221 8128 4229 8192
rect 3909 8127 4229 8128
rect 9840 8192 10160 8193
rect 9840 8128 9848 8192
rect 9912 8128 9928 8192
rect 9992 8128 10008 8192
rect 10072 8128 10088 8192
rect 10152 8128 10160 8192
rect 9840 8127 10160 8128
rect 15770 8192 16090 8193
rect 15770 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15938 8192
rect 16002 8128 16018 8192
rect 16082 8128 16090 8192
rect 15770 8127 16090 8128
rect 6874 7648 7194 7649
rect 6874 7584 6882 7648
rect 6946 7584 6962 7648
rect 7026 7584 7042 7648
rect 7106 7584 7122 7648
rect 7186 7584 7194 7648
rect 6874 7583 7194 7584
rect 12805 7648 13125 7649
rect 12805 7584 12813 7648
rect 12877 7584 12893 7648
rect 12957 7584 12973 7648
rect 13037 7584 13053 7648
rect 13117 7584 13125 7648
rect 12805 7583 13125 7584
rect 3909 7104 4229 7105
rect 3909 7040 3917 7104
rect 3981 7040 3997 7104
rect 4061 7040 4077 7104
rect 4141 7040 4157 7104
rect 4221 7040 4229 7104
rect 3909 7039 4229 7040
rect 9840 7104 10160 7105
rect 9840 7040 9848 7104
rect 9912 7040 9928 7104
rect 9992 7040 10008 7104
rect 10072 7040 10088 7104
rect 10152 7040 10160 7104
rect 9840 7039 10160 7040
rect 15770 7104 16090 7105
rect 15770 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15938 7104
rect 16002 7040 16018 7104
rect 16082 7040 16090 7104
rect 15770 7039 16090 7040
rect 6874 6560 7194 6561
rect 6874 6496 6882 6560
rect 6946 6496 6962 6560
rect 7026 6496 7042 6560
rect 7106 6496 7122 6560
rect 7186 6496 7194 6560
rect 6874 6495 7194 6496
rect 12805 6560 13125 6561
rect 12805 6496 12813 6560
rect 12877 6496 12893 6560
rect 12957 6496 12973 6560
rect 13037 6496 13053 6560
rect 13117 6496 13125 6560
rect 12805 6495 13125 6496
rect 3909 6016 4229 6017
rect 3909 5952 3917 6016
rect 3981 5952 3997 6016
rect 4061 5952 4077 6016
rect 4141 5952 4157 6016
rect 4221 5952 4229 6016
rect 3909 5951 4229 5952
rect 9840 6016 10160 6017
rect 9840 5952 9848 6016
rect 9912 5952 9928 6016
rect 9992 5952 10008 6016
rect 10072 5952 10088 6016
rect 10152 5952 10160 6016
rect 9840 5951 10160 5952
rect 15770 6016 16090 6017
rect 15770 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15938 6016
rect 16002 5952 16018 6016
rect 16082 5952 16090 6016
rect 15770 5951 16090 5952
rect 6874 5472 7194 5473
rect 6874 5408 6882 5472
rect 6946 5408 6962 5472
rect 7026 5408 7042 5472
rect 7106 5408 7122 5472
rect 7186 5408 7194 5472
rect 6874 5407 7194 5408
rect 12805 5472 13125 5473
rect 12805 5408 12813 5472
rect 12877 5408 12893 5472
rect 12957 5408 12973 5472
rect 13037 5408 13053 5472
rect 13117 5408 13125 5472
rect 12805 5407 13125 5408
rect 3909 4928 4229 4929
rect 3909 4864 3917 4928
rect 3981 4864 3997 4928
rect 4061 4864 4077 4928
rect 4141 4864 4157 4928
rect 4221 4864 4229 4928
rect 3909 4863 4229 4864
rect 9840 4928 10160 4929
rect 9840 4864 9848 4928
rect 9912 4864 9928 4928
rect 9992 4864 10008 4928
rect 10072 4864 10088 4928
rect 10152 4864 10160 4928
rect 9840 4863 10160 4864
rect 15770 4928 16090 4929
rect 15770 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15938 4928
rect 16002 4864 16018 4928
rect 16082 4864 16090 4928
rect 15770 4863 16090 4864
rect 6874 4384 7194 4385
rect 6874 4320 6882 4384
rect 6946 4320 6962 4384
rect 7026 4320 7042 4384
rect 7106 4320 7122 4384
rect 7186 4320 7194 4384
rect 6874 4319 7194 4320
rect 12805 4384 13125 4385
rect 12805 4320 12813 4384
rect 12877 4320 12893 4384
rect 12957 4320 12973 4384
rect 13037 4320 13053 4384
rect 13117 4320 13125 4384
rect 12805 4319 13125 4320
rect 3909 3840 4229 3841
rect 3909 3776 3917 3840
rect 3981 3776 3997 3840
rect 4061 3776 4077 3840
rect 4141 3776 4157 3840
rect 4221 3776 4229 3840
rect 3909 3775 4229 3776
rect 9840 3840 10160 3841
rect 9840 3776 9848 3840
rect 9912 3776 9928 3840
rect 9992 3776 10008 3840
rect 10072 3776 10088 3840
rect 10152 3776 10160 3840
rect 9840 3775 10160 3776
rect 15770 3840 16090 3841
rect 15770 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15938 3840
rect 16002 3776 16018 3840
rect 16082 3776 16090 3840
rect 15770 3775 16090 3776
rect 6874 3296 7194 3297
rect 6874 3232 6882 3296
rect 6946 3232 6962 3296
rect 7026 3232 7042 3296
rect 7106 3232 7122 3296
rect 7186 3232 7194 3296
rect 6874 3231 7194 3232
rect 12805 3296 13125 3297
rect 12805 3232 12813 3296
rect 12877 3232 12893 3296
rect 12957 3232 12973 3296
rect 13037 3232 13053 3296
rect 13117 3232 13125 3296
rect 12805 3231 13125 3232
rect 18045 3226 18111 3229
rect 19200 3226 20000 3256
rect 18045 3224 20000 3226
rect 18045 3168 18050 3224
rect 18106 3168 20000 3224
rect 18045 3166 20000 3168
rect 18045 3163 18111 3166
rect 19200 3136 20000 3166
rect 2221 2954 2287 2957
rect 16614 2954 16620 2956
rect 2221 2952 16620 2954
rect 2221 2896 2226 2952
rect 2282 2896 16620 2952
rect 2221 2894 16620 2896
rect 2221 2891 2287 2894
rect 16614 2892 16620 2894
rect 16684 2892 16690 2956
rect 0 2818 800 2848
rect 1485 2818 1551 2821
rect 0 2816 1551 2818
rect 0 2760 1490 2816
rect 1546 2760 1551 2816
rect 0 2758 1551 2760
rect 0 2728 800 2758
rect 1485 2755 1551 2758
rect 3909 2752 4229 2753
rect 3909 2688 3917 2752
rect 3981 2688 3997 2752
rect 4061 2688 4077 2752
rect 4141 2688 4157 2752
rect 4221 2688 4229 2752
rect 3909 2687 4229 2688
rect 9840 2752 10160 2753
rect 9840 2688 9848 2752
rect 9912 2688 9928 2752
rect 9992 2688 10008 2752
rect 10072 2688 10088 2752
rect 10152 2688 10160 2752
rect 9840 2687 10160 2688
rect 15770 2752 16090 2753
rect 15770 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15938 2752
rect 16002 2688 16018 2752
rect 16082 2688 16090 2752
rect 15770 2687 16090 2688
rect 6874 2208 7194 2209
rect 6874 2144 6882 2208
rect 6946 2144 6962 2208
rect 7026 2144 7042 2208
rect 7106 2144 7122 2208
rect 7186 2144 7194 2208
rect 6874 2143 7194 2144
rect 12805 2208 13125 2209
rect 12805 2144 12813 2208
rect 12877 2144 12893 2208
rect 12957 2144 12973 2208
rect 13037 2144 13053 2208
rect 13117 2144 13125 2208
rect 12805 2143 13125 2144
<< via3 >>
rect 3917 47356 3981 47360
rect 3917 47300 3921 47356
rect 3921 47300 3977 47356
rect 3977 47300 3981 47356
rect 3917 47296 3981 47300
rect 3997 47356 4061 47360
rect 3997 47300 4001 47356
rect 4001 47300 4057 47356
rect 4057 47300 4061 47356
rect 3997 47296 4061 47300
rect 4077 47356 4141 47360
rect 4077 47300 4081 47356
rect 4081 47300 4137 47356
rect 4137 47300 4141 47356
rect 4077 47296 4141 47300
rect 4157 47356 4221 47360
rect 4157 47300 4161 47356
rect 4161 47300 4217 47356
rect 4217 47300 4221 47356
rect 4157 47296 4221 47300
rect 9848 47356 9912 47360
rect 9848 47300 9852 47356
rect 9852 47300 9908 47356
rect 9908 47300 9912 47356
rect 9848 47296 9912 47300
rect 9928 47356 9992 47360
rect 9928 47300 9932 47356
rect 9932 47300 9988 47356
rect 9988 47300 9992 47356
rect 9928 47296 9992 47300
rect 10008 47356 10072 47360
rect 10008 47300 10012 47356
rect 10012 47300 10068 47356
rect 10068 47300 10072 47356
rect 10008 47296 10072 47300
rect 10088 47356 10152 47360
rect 10088 47300 10092 47356
rect 10092 47300 10148 47356
rect 10148 47300 10152 47356
rect 10088 47296 10152 47300
rect 15778 47356 15842 47360
rect 15778 47300 15782 47356
rect 15782 47300 15838 47356
rect 15838 47300 15842 47356
rect 15778 47296 15842 47300
rect 15858 47356 15922 47360
rect 15858 47300 15862 47356
rect 15862 47300 15918 47356
rect 15918 47300 15922 47356
rect 15858 47296 15922 47300
rect 15938 47356 16002 47360
rect 15938 47300 15942 47356
rect 15942 47300 15998 47356
rect 15998 47300 16002 47356
rect 15938 47296 16002 47300
rect 16018 47356 16082 47360
rect 16018 47300 16022 47356
rect 16022 47300 16078 47356
rect 16078 47300 16082 47356
rect 16018 47296 16082 47300
rect 6882 46812 6946 46816
rect 6882 46756 6886 46812
rect 6886 46756 6942 46812
rect 6942 46756 6946 46812
rect 6882 46752 6946 46756
rect 6962 46812 7026 46816
rect 6962 46756 6966 46812
rect 6966 46756 7022 46812
rect 7022 46756 7026 46812
rect 6962 46752 7026 46756
rect 7042 46812 7106 46816
rect 7042 46756 7046 46812
rect 7046 46756 7102 46812
rect 7102 46756 7106 46812
rect 7042 46752 7106 46756
rect 7122 46812 7186 46816
rect 7122 46756 7126 46812
rect 7126 46756 7182 46812
rect 7182 46756 7186 46812
rect 7122 46752 7186 46756
rect 12813 46812 12877 46816
rect 12813 46756 12817 46812
rect 12817 46756 12873 46812
rect 12873 46756 12877 46812
rect 12813 46752 12877 46756
rect 12893 46812 12957 46816
rect 12893 46756 12897 46812
rect 12897 46756 12953 46812
rect 12953 46756 12957 46812
rect 12893 46752 12957 46756
rect 12973 46812 13037 46816
rect 12973 46756 12977 46812
rect 12977 46756 13033 46812
rect 13033 46756 13037 46812
rect 12973 46752 13037 46756
rect 13053 46812 13117 46816
rect 13053 46756 13057 46812
rect 13057 46756 13113 46812
rect 13113 46756 13117 46812
rect 13053 46752 13117 46756
rect 3917 46268 3981 46272
rect 3917 46212 3921 46268
rect 3921 46212 3977 46268
rect 3977 46212 3981 46268
rect 3917 46208 3981 46212
rect 3997 46268 4061 46272
rect 3997 46212 4001 46268
rect 4001 46212 4057 46268
rect 4057 46212 4061 46268
rect 3997 46208 4061 46212
rect 4077 46268 4141 46272
rect 4077 46212 4081 46268
rect 4081 46212 4137 46268
rect 4137 46212 4141 46268
rect 4077 46208 4141 46212
rect 4157 46268 4221 46272
rect 4157 46212 4161 46268
rect 4161 46212 4217 46268
rect 4217 46212 4221 46268
rect 4157 46208 4221 46212
rect 9848 46268 9912 46272
rect 9848 46212 9852 46268
rect 9852 46212 9908 46268
rect 9908 46212 9912 46268
rect 9848 46208 9912 46212
rect 9928 46268 9992 46272
rect 9928 46212 9932 46268
rect 9932 46212 9988 46268
rect 9988 46212 9992 46268
rect 9928 46208 9992 46212
rect 10008 46268 10072 46272
rect 10008 46212 10012 46268
rect 10012 46212 10068 46268
rect 10068 46212 10072 46268
rect 10008 46208 10072 46212
rect 10088 46268 10152 46272
rect 10088 46212 10092 46268
rect 10092 46212 10148 46268
rect 10148 46212 10152 46268
rect 10088 46208 10152 46212
rect 15778 46268 15842 46272
rect 15778 46212 15782 46268
rect 15782 46212 15838 46268
rect 15838 46212 15842 46268
rect 15778 46208 15842 46212
rect 15858 46268 15922 46272
rect 15858 46212 15862 46268
rect 15862 46212 15918 46268
rect 15918 46212 15922 46268
rect 15858 46208 15922 46212
rect 15938 46268 16002 46272
rect 15938 46212 15942 46268
rect 15942 46212 15998 46268
rect 15998 46212 16002 46268
rect 15938 46208 16002 46212
rect 16018 46268 16082 46272
rect 16018 46212 16022 46268
rect 16022 46212 16078 46268
rect 16078 46212 16082 46268
rect 16018 46208 16082 46212
rect 15516 45928 15580 45932
rect 15516 45872 15566 45928
rect 15566 45872 15580 45928
rect 15516 45868 15580 45872
rect 6882 45724 6946 45728
rect 6882 45668 6886 45724
rect 6886 45668 6942 45724
rect 6942 45668 6946 45724
rect 6882 45664 6946 45668
rect 6962 45724 7026 45728
rect 6962 45668 6966 45724
rect 6966 45668 7022 45724
rect 7022 45668 7026 45724
rect 6962 45664 7026 45668
rect 7042 45724 7106 45728
rect 7042 45668 7046 45724
rect 7046 45668 7102 45724
rect 7102 45668 7106 45724
rect 7042 45664 7106 45668
rect 7122 45724 7186 45728
rect 7122 45668 7126 45724
rect 7126 45668 7182 45724
rect 7182 45668 7186 45724
rect 7122 45664 7186 45668
rect 12813 45724 12877 45728
rect 12813 45668 12817 45724
rect 12817 45668 12873 45724
rect 12873 45668 12877 45724
rect 12813 45664 12877 45668
rect 12893 45724 12957 45728
rect 12893 45668 12897 45724
rect 12897 45668 12953 45724
rect 12953 45668 12957 45724
rect 12893 45664 12957 45668
rect 12973 45724 13037 45728
rect 12973 45668 12977 45724
rect 12977 45668 13033 45724
rect 13033 45668 13037 45724
rect 12973 45664 13037 45668
rect 13053 45724 13117 45728
rect 13053 45668 13057 45724
rect 13057 45668 13113 45724
rect 13113 45668 13117 45724
rect 13053 45664 13117 45668
rect 3917 45180 3981 45184
rect 3917 45124 3921 45180
rect 3921 45124 3977 45180
rect 3977 45124 3981 45180
rect 3917 45120 3981 45124
rect 3997 45180 4061 45184
rect 3997 45124 4001 45180
rect 4001 45124 4057 45180
rect 4057 45124 4061 45180
rect 3997 45120 4061 45124
rect 4077 45180 4141 45184
rect 4077 45124 4081 45180
rect 4081 45124 4137 45180
rect 4137 45124 4141 45180
rect 4077 45120 4141 45124
rect 4157 45180 4221 45184
rect 4157 45124 4161 45180
rect 4161 45124 4217 45180
rect 4217 45124 4221 45180
rect 4157 45120 4221 45124
rect 9848 45180 9912 45184
rect 9848 45124 9852 45180
rect 9852 45124 9908 45180
rect 9908 45124 9912 45180
rect 9848 45120 9912 45124
rect 9928 45180 9992 45184
rect 9928 45124 9932 45180
rect 9932 45124 9988 45180
rect 9988 45124 9992 45180
rect 9928 45120 9992 45124
rect 10008 45180 10072 45184
rect 10008 45124 10012 45180
rect 10012 45124 10068 45180
rect 10068 45124 10072 45180
rect 10008 45120 10072 45124
rect 10088 45180 10152 45184
rect 10088 45124 10092 45180
rect 10092 45124 10148 45180
rect 10148 45124 10152 45180
rect 10088 45120 10152 45124
rect 15778 45180 15842 45184
rect 15778 45124 15782 45180
rect 15782 45124 15838 45180
rect 15838 45124 15842 45180
rect 15778 45120 15842 45124
rect 15858 45180 15922 45184
rect 15858 45124 15862 45180
rect 15862 45124 15918 45180
rect 15918 45124 15922 45180
rect 15858 45120 15922 45124
rect 15938 45180 16002 45184
rect 15938 45124 15942 45180
rect 15942 45124 15998 45180
rect 15998 45124 16002 45180
rect 15938 45120 16002 45124
rect 16018 45180 16082 45184
rect 16018 45124 16022 45180
rect 16022 45124 16078 45180
rect 16078 45124 16082 45180
rect 16018 45120 16082 45124
rect 6882 44636 6946 44640
rect 6882 44580 6886 44636
rect 6886 44580 6942 44636
rect 6942 44580 6946 44636
rect 6882 44576 6946 44580
rect 6962 44636 7026 44640
rect 6962 44580 6966 44636
rect 6966 44580 7022 44636
rect 7022 44580 7026 44636
rect 6962 44576 7026 44580
rect 7042 44636 7106 44640
rect 7042 44580 7046 44636
rect 7046 44580 7102 44636
rect 7102 44580 7106 44636
rect 7042 44576 7106 44580
rect 7122 44636 7186 44640
rect 7122 44580 7126 44636
rect 7126 44580 7182 44636
rect 7182 44580 7186 44636
rect 7122 44576 7186 44580
rect 12813 44636 12877 44640
rect 12813 44580 12817 44636
rect 12817 44580 12873 44636
rect 12873 44580 12877 44636
rect 12813 44576 12877 44580
rect 12893 44636 12957 44640
rect 12893 44580 12897 44636
rect 12897 44580 12953 44636
rect 12953 44580 12957 44636
rect 12893 44576 12957 44580
rect 12973 44636 13037 44640
rect 12973 44580 12977 44636
rect 12977 44580 13033 44636
rect 13033 44580 13037 44636
rect 12973 44576 13037 44580
rect 13053 44636 13117 44640
rect 13053 44580 13057 44636
rect 13057 44580 13113 44636
rect 13113 44580 13117 44636
rect 13053 44576 13117 44580
rect 3917 44092 3981 44096
rect 3917 44036 3921 44092
rect 3921 44036 3977 44092
rect 3977 44036 3981 44092
rect 3917 44032 3981 44036
rect 3997 44092 4061 44096
rect 3997 44036 4001 44092
rect 4001 44036 4057 44092
rect 4057 44036 4061 44092
rect 3997 44032 4061 44036
rect 4077 44092 4141 44096
rect 4077 44036 4081 44092
rect 4081 44036 4137 44092
rect 4137 44036 4141 44092
rect 4077 44032 4141 44036
rect 4157 44092 4221 44096
rect 4157 44036 4161 44092
rect 4161 44036 4217 44092
rect 4217 44036 4221 44092
rect 4157 44032 4221 44036
rect 9848 44092 9912 44096
rect 9848 44036 9852 44092
rect 9852 44036 9908 44092
rect 9908 44036 9912 44092
rect 9848 44032 9912 44036
rect 9928 44092 9992 44096
rect 9928 44036 9932 44092
rect 9932 44036 9988 44092
rect 9988 44036 9992 44092
rect 9928 44032 9992 44036
rect 10008 44092 10072 44096
rect 10008 44036 10012 44092
rect 10012 44036 10068 44092
rect 10068 44036 10072 44092
rect 10008 44032 10072 44036
rect 10088 44092 10152 44096
rect 10088 44036 10092 44092
rect 10092 44036 10148 44092
rect 10148 44036 10152 44092
rect 10088 44032 10152 44036
rect 15778 44092 15842 44096
rect 15778 44036 15782 44092
rect 15782 44036 15838 44092
rect 15838 44036 15842 44092
rect 15778 44032 15842 44036
rect 15858 44092 15922 44096
rect 15858 44036 15862 44092
rect 15862 44036 15918 44092
rect 15918 44036 15922 44092
rect 15858 44032 15922 44036
rect 15938 44092 16002 44096
rect 15938 44036 15942 44092
rect 15942 44036 15998 44092
rect 15998 44036 16002 44092
rect 15938 44032 16002 44036
rect 16018 44092 16082 44096
rect 16018 44036 16022 44092
rect 16022 44036 16078 44092
rect 16078 44036 16082 44092
rect 16018 44032 16082 44036
rect 6882 43548 6946 43552
rect 6882 43492 6886 43548
rect 6886 43492 6942 43548
rect 6942 43492 6946 43548
rect 6882 43488 6946 43492
rect 6962 43548 7026 43552
rect 6962 43492 6966 43548
rect 6966 43492 7022 43548
rect 7022 43492 7026 43548
rect 6962 43488 7026 43492
rect 7042 43548 7106 43552
rect 7042 43492 7046 43548
rect 7046 43492 7102 43548
rect 7102 43492 7106 43548
rect 7042 43488 7106 43492
rect 7122 43548 7186 43552
rect 7122 43492 7126 43548
rect 7126 43492 7182 43548
rect 7182 43492 7186 43548
rect 7122 43488 7186 43492
rect 12813 43548 12877 43552
rect 12813 43492 12817 43548
rect 12817 43492 12873 43548
rect 12873 43492 12877 43548
rect 12813 43488 12877 43492
rect 12893 43548 12957 43552
rect 12893 43492 12897 43548
rect 12897 43492 12953 43548
rect 12953 43492 12957 43548
rect 12893 43488 12957 43492
rect 12973 43548 13037 43552
rect 12973 43492 12977 43548
rect 12977 43492 13033 43548
rect 13033 43492 13037 43548
rect 12973 43488 13037 43492
rect 13053 43548 13117 43552
rect 13053 43492 13057 43548
rect 13057 43492 13113 43548
rect 13113 43492 13117 43548
rect 13053 43488 13117 43492
rect 3917 43004 3981 43008
rect 3917 42948 3921 43004
rect 3921 42948 3977 43004
rect 3977 42948 3981 43004
rect 3917 42944 3981 42948
rect 3997 43004 4061 43008
rect 3997 42948 4001 43004
rect 4001 42948 4057 43004
rect 4057 42948 4061 43004
rect 3997 42944 4061 42948
rect 4077 43004 4141 43008
rect 4077 42948 4081 43004
rect 4081 42948 4137 43004
rect 4137 42948 4141 43004
rect 4077 42944 4141 42948
rect 4157 43004 4221 43008
rect 4157 42948 4161 43004
rect 4161 42948 4217 43004
rect 4217 42948 4221 43004
rect 4157 42944 4221 42948
rect 9848 43004 9912 43008
rect 9848 42948 9852 43004
rect 9852 42948 9908 43004
rect 9908 42948 9912 43004
rect 9848 42944 9912 42948
rect 9928 43004 9992 43008
rect 9928 42948 9932 43004
rect 9932 42948 9988 43004
rect 9988 42948 9992 43004
rect 9928 42944 9992 42948
rect 10008 43004 10072 43008
rect 10008 42948 10012 43004
rect 10012 42948 10068 43004
rect 10068 42948 10072 43004
rect 10008 42944 10072 42948
rect 10088 43004 10152 43008
rect 10088 42948 10092 43004
rect 10092 42948 10148 43004
rect 10148 42948 10152 43004
rect 10088 42944 10152 42948
rect 15778 43004 15842 43008
rect 15778 42948 15782 43004
rect 15782 42948 15838 43004
rect 15838 42948 15842 43004
rect 15778 42944 15842 42948
rect 15858 43004 15922 43008
rect 15858 42948 15862 43004
rect 15862 42948 15918 43004
rect 15918 42948 15922 43004
rect 15858 42944 15922 42948
rect 15938 43004 16002 43008
rect 15938 42948 15942 43004
rect 15942 42948 15998 43004
rect 15998 42948 16002 43004
rect 15938 42944 16002 42948
rect 16018 43004 16082 43008
rect 16018 42948 16022 43004
rect 16022 42948 16078 43004
rect 16078 42948 16082 43004
rect 16018 42944 16082 42948
rect 6882 42460 6946 42464
rect 6882 42404 6886 42460
rect 6886 42404 6942 42460
rect 6942 42404 6946 42460
rect 6882 42400 6946 42404
rect 6962 42460 7026 42464
rect 6962 42404 6966 42460
rect 6966 42404 7022 42460
rect 7022 42404 7026 42460
rect 6962 42400 7026 42404
rect 7042 42460 7106 42464
rect 7042 42404 7046 42460
rect 7046 42404 7102 42460
rect 7102 42404 7106 42460
rect 7042 42400 7106 42404
rect 7122 42460 7186 42464
rect 7122 42404 7126 42460
rect 7126 42404 7182 42460
rect 7182 42404 7186 42460
rect 7122 42400 7186 42404
rect 12813 42460 12877 42464
rect 12813 42404 12817 42460
rect 12817 42404 12873 42460
rect 12873 42404 12877 42460
rect 12813 42400 12877 42404
rect 12893 42460 12957 42464
rect 12893 42404 12897 42460
rect 12897 42404 12953 42460
rect 12953 42404 12957 42460
rect 12893 42400 12957 42404
rect 12973 42460 13037 42464
rect 12973 42404 12977 42460
rect 12977 42404 13033 42460
rect 13033 42404 13037 42460
rect 12973 42400 13037 42404
rect 13053 42460 13117 42464
rect 13053 42404 13057 42460
rect 13057 42404 13113 42460
rect 13113 42404 13117 42460
rect 13053 42400 13117 42404
rect 3917 41916 3981 41920
rect 3917 41860 3921 41916
rect 3921 41860 3977 41916
rect 3977 41860 3981 41916
rect 3917 41856 3981 41860
rect 3997 41916 4061 41920
rect 3997 41860 4001 41916
rect 4001 41860 4057 41916
rect 4057 41860 4061 41916
rect 3997 41856 4061 41860
rect 4077 41916 4141 41920
rect 4077 41860 4081 41916
rect 4081 41860 4137 41916
rect 4137 41860 4141 41916
rect 4077 41856 4141 41860
rect 4157 41916 4221 41920
rect 4157 41860 4161 41916
rect 4161 41860 4217 41916
rect 4217 41860 4221 41916
rect 4157 41856 4221 41860
rect 9848 41916 9912 41920
rect 9848 41860 9852 41916
rect 9852 41860 9908 41916
rect 9908 41860 9912 41916
rect 9848 41856 9912 41860
rect 9928 41916 9992 41920
rect 9928 41860 9932 41916
rect 9932 41860 9988 41916
rect 9988 41860 9992 41916
rect 9928 41856 9992 41860
rect 10008 41916 10072 41920
rect 10008 41860 10012 41916
rect 10012 41860 10068 41916
rect 10068 41860 10072 41916
rect 10008 41856 10072 41860
rect 10088 41916 10152 41920
rect 10088 41860 10092 41916
rect 10092 41860 10148 41916
rect 10148 41860 10152 41916
rect 10088 41856 10152 41860
rect 15778 41916 15842 41920
rect 15778 41860 15782 41916
rect 15782 41860 15838 41916
rect 15838 41860 15842 41916
rect 15778 41856 15842 41860
rect 15858 41916 15922 41920
rect 15858 41860 15862 41916
rect 15862 41860 15918 41916
rect 15918 41860 15922 41916
rect 15858 41856 15922 41860
rect 15938 41916 16002 41920
rect 15938 41860 15942 41916
rect 15942 41860 15998 41916
rect 15998 41860 16002 41916
rect 15938 41856 16002 41860
rect 16018 41916 16082 41920
rect 16018 41860 16022 41916
rect 16022 41860 16078 41916
rect 16078 41860 16082 41916
rect 16018 41856 16082 41860
rect 6882 41372 6946 41376
rect 6882 41316 6886 41372
rect 6886 41316 6942 41372
rect 6942 41316 6946 41372
rect 6882 41312 6946 41316
rect 6962 41372 7026 41376
rect 6962 41316 6966 41372
rect 6966 41316 7022 41372
rect 7022 41316 7026 41372
rect 6962 41312 7026 41316
rect 7042 41372 7106 41376
rect 7042 41316 7046 41372
rect 7046 41316 7102 41372
rect 7102 41316 7106 41372
rect 7042 41312 7106 41316
rect 7122 41372 7186 41376
rect 7122 41316 7126 41372
rect 7126 41316 7182 41372
rect 7182 41316 7186 41372
rect 7122 41312 7186 41316
rect 12813 41372 12877 41376
rect 12813 41316 12817 41372
rect 12817 41316 12873 41372
rect 12873 41316 12877 41372
rect 12813 41312 12877 41316
rect 12893 41372 12957 41376
rect 12893 41316 12897 41372
rect 12897 41316 12953 41372
rect 12953 41316 12957 41372
rect 12893 41312 12957 41316
rect 12973 41372 13037 41376
rect 12973 41316 12977 41372
rect 12977 41316 13033 41372
rect 13033 41316 13037 41372
rect 12973 41312 13037 41316
rect 13053 41372 13117 41376
rect 13053 41316 13057 41372
rect 13057 41316 13113 41372
rect 13113 41316 13117 41372
rect 13053 41312 13117 41316
rect 3917 40828 3981 40832
rect 3917 40772 3921 40828
rect 3921 40772 3977 40828
rect 3977 40772 3981 40828
rect 3917 40768 3981 40772
rect 3997 40828 4061 40832
rect 3997 40772 4001 40828
rect 4001 40772 4057 40828
rect 4057 40772 4061 40828
rect 3997 40768 4061 40772
rect 4077 40828 4141 40832
rect 4077 40772 4081 40828
rect 4081 40772 4137 40828
rect 4137 40772 4141 40828
rect 4077 40768 4141 40772
rect 4157 40828 4221 40832
rect 4157 40772 4161 40828
rect 4161 40772 4217 40828
rect 4217 40772 4221 40828
rect 4157 40768 4221 40772
rect 9848 40828 9912 40832
rect 9848 40772 9852 40828
rect 9852 40772 9908 40828
rect 9908 40772 9912 40828
rect 9848 40768 9912 40772
rect 9928 40828 9992 40832
rect 9928 40772 9932 40828
rect 9932 40772 9988 40828
rect 9988 40772 9992 40828
rect 9928 40768 9992 40772
rect 10008 40828 10072 40832
rect 10008 40772 10012 40828
rect 10012 40772 10068 40828
rect 10068 40772 10072 40828
rect 10008 40768 10072 40772
rect 10088 40828 10152 40832
rect 10088 40772 10092 40828
rect 10092 40772 10148 40828
rect 10148 40772 10152 40828
rect 10088 40768 10152 40772
rect 15778 40828 15842 40832
rect 15778 40772 15782 40828
rect 15782 40772 15838 40828
rect 15838 40772 15842 40828
rect 15778 40768 15842 40772
rect 15858 40828 15922 40832
rect 15858 40772 15862 40828
rect 15862 40772 15918 40828
rect 15918 40772 15922 40828
rect 15858 40768 15922 40772
rect 15938 40828 16002 40832
rect 15938 40772 15942 40828
rect 15942 40772 15998 40828
rect 15998 40772 16002 40828
rect 15938 40768 16002 40772
rect 16018 40828 16082 40832
rect 16018 40772 16022 40828
rect 16022 40772 16078 40828
rect 16078 40772 16082 40828
rect 16018 40768 16082 40772
rect 6882 40284 6946 40288
rect 6882 40228 6886 40284
rect 6886 40228 6942 40284
rect 6942 40228 6946 40284
rect 6882 40224 6946 40228
rect 6962 40284 7026 40288
rect 6962 40228 6966 40284
rect 6966 40228 7022 40284
rect 7022 40228 7026 40284
rect 6962 40224 7026 40228
rect 7042 40284 7106 40288
rect 7042 40228 7046 40284
rect 7046 40228 7102 40284
rect 7102 40228 7106 40284
rect 7042 40224 7106 40228
rect 7122 40284 7186 40288
rect 7122 40228 7126 40284
rect 7126 40228 7182 40284
rect 7182 40228 7186 40284
rect 7122 40224 7186 40228
rect 12813 40284 12877 40288
rect 12813 40228 12817 40284
rect 12817 40228 12873 40284
rect 12873 40228 12877 40284
rect 12813 40224 12877 40228
rect 12893 40284 12957 40288
rect 12893 40228 12897 40284
rect 12897 40228 12953 40284
rect 12953 40228 12957 40284
rect 12893 40224 12957 40228
rect 12973 40284 13037 40288
rect 12973 40228 12977 40284
rect 12977 40228 13033 40284
rect 13033 40228 13037 40284
rect 12973 40224 13037 40228
rect 13053 40284 13117 40288
rect 13053 40228 13057 40284
rect 13057 40228 13113 40284
rect 13113 40228 13117 40284
rect 13053 40224 13117 40228
rect 3917 39740 3981 39744
rect 3917 39684 3921 39740
rect 3921 39684 3977 39740
rect 3977 39684 3981 39740
rect 3917 39680 3981 39684
rect 3997 39740 4061 39744
rect 3997 39684 4001 39740
rect 4001 39684 4057 39740
rect 4057 39684 4061 39740
rect 3997 39680 4061 39684
rect 4077 39740 4141 39744
rect 4077 39684 4081 39740
rect 4081 39684 4137 39740
rect 4137 39684 4141 39740
rect 4077 39680 4141 39684
rect 4157 39740 4221 39744
rect 4157 39684 4161 39740
rect 4161 39684 4217 39740
rect 4217 39684 4221 39740
rect 4157 39680 4221 39684
rect 9848 39740 9912 39744
rect 9848 39684 9852 39740
rect 9852 39684 9908 39740
rect 9908 39684 9912 39740
rect 9848 39680 9912 39684
rect 9928 39740 9992 39744
rect 9928 39684 9932 39740
rect 9932 39684 9988 39740
rect 9988 39684 9992 39740
rect 9928 39680 9992 39684
rect 10008 39740 10072 39744
rect 10008 39684 10012 39740
rect 10012 39684 10068 39740
rect 10068 39684 10072 39740
rect 10008 39680 10072 39684
rect 10088 39740 10152 39744
rect 10088 39684 10092 39740
rect 10092 39684 10148 39740
rect 10148 39684 10152 39740
rect 10088 39680 10152 39684
rect 15778 39740 15842 39744
rect 15778 39684 15782 39740
rect 15782 39684 15838 39740
rect 15838 39684 15842 39740
rect 15778 39680 15842 39684
rect 15858 39740 15922 39744
rect 15858 39684 15862 39740
rect 15862 39684 15918 39740
rect 15918 39684 15922 39740
rect 15858 39680 15922 39684
rect 15938 39740 16002 39744
rect 15938 39684 15942 39740
rect 15942 39684 15998 39740
rect 15998 39684 16002 39740
rect 15938 39680 16002 39684
rect 16018 39740 16082 39744
rect 16018 39684 16022 39740
rect 16022 39684 16078 39740
rect 16078 39684 16082 39740
rect 16018 39680 16082 39684
rect 6882 39196 6946 39200
rect 6882 39140 6886 39196
rect 6886 39140 6942 39196
rect 6942 39140 6946 39196
rect 6882 39136 6946 39140
rect 6962 39196 7026 39200
rect 6962 39140 6966 39196
rect 6966 39140 7022 39196
rect 7022 39140 7026 39196
rect 6962 39136 7026 39140
rect 7042 39196 7106 39200
rect 7042 39140 7046 39196
rect 7046 39140 7102 39196
rect 7102 39140 7106 39196
rect 7042 39136 7106 39140
rect 7122 39196 7186 39200
rect 7122 39140 7126 39196
rect 7126 39140 7182 39196
rect 7182 39140 7186 39196
rect 7122 39136 7186 39140
rect 12813 39196 12877 39200
rect 12813 39140 12817 39196
rect 12817 39140 12873 39196
rect 12873 39140 12877 39196
rect 12813 39136 12877 39140
rect 12893 39196 12957 39200
rect 12893 39140 12897 39196
rect 12897 39140 12953 39196
rect 12953 39140 12957 39196
rect 12893 39136 12957 39140
rect 12973 39196 13037 39200
rect 12973 39140 12977 39196
rect 12977 39140 13033 39196
rect 13033 39140 13037 39196
rect 12973 39136 13037 39140
rect 13053 39196 13117 39200
rect 13053 39140 13057 39196
rect 13057 39140 13113 39196
rect 13113 39140 13117 39196
rect 13053 39136 13117 39140
rect 3917 38652 3981 38656
rect 3917 38596 3921 38652
rect 3921 38596 3977 38652
rect 3977 38596 3981 38652
rect 3917 38592 3981 38596
rect 3997 38652 4061 38656
rect 3997 38596 4001 38652
rect 4001 38596 4057 38652
rect 4057 38596 4061 38652
rect 3997 38592 4061 38596
rect 4077 38652 4141 38656
rect 4077 38596 4081 38652
rect 4081 38596 4137 38652
rect 4137 38596 4141 38652
rect 4077 38592 4141 38596
rect 4157 38652 4221 38656
rect 4157 38596 4161 38652
rect 4161 38596 4217 38652
rect 4217 38596 4221 38652
rect 4157 38592 4221 38596
rect 9848 38652 9912 38656
rect 9848 38596 9852 38652
rect 9852 38596 9908 38652
rect 9908 38596 9912 38652
rect 9848 38592 9912 38596
rect 9928 38652 9992 38656
rect 9928 38596 9932 38652
rect 9932 38596 9988 38652
rect 9988 38596 9992 38652
rect 9928 38592 9992 38596
rect 10008 38652 10072 38656
rect 10008 38596 10012 38652
rect 10012 38596 10068 38652
rect 10068 38596 10072 38652
rect 10008 38592 10072 38596
rect 10088 38652 10152 38656
rect 10088 38596 10092 38652
rect 10092 38596 10148 38652
rect 10148 38596 10152 38652
rect 10088 38592 10152 38596
rect 15778 38652 15842 38656
rect 15778 38596 15782 38652
rect 15782 38596 15838 38652
rect 15838 38596 15842 38652
rect 15778 38592 15842 38596
rect 15858 38652 15922 38656
rect 15858 38596 15862 38652
rect 15862 38596 15918 38652
rect 15918 38596 15922 38652
rect 15858 38592 15922 38596
rect 15938 38652 16002 38656
rect 15938 38596 15942 38652
rect 15942 38596 15998 38652
rect 15998 38596 16002 38652
rect 15938 38592 16002 38596
rect 16018 38652 16082 38656
rect 16018 38596 16022 38652
rect 16022 38596 16078 38652
rect 16078 38596 16082 38652
rect 16018 38592 16082 38596
rect 6882 38108 6946 38112
rect 6882 38052 6886 38108
rect 6886 38052 6942 38108
rect 6942 38052 6946 38108
rect 6882 38048 6946 38052
rect 6962 38108 7026 38112
rect 6962 38052 6966 38108
rect 6966 38052 7022 38108
rect 7022 38052 7026 38108
rect 6962 38048 7026 38052
rect 7042 38108 7106 38112
rect 7042 38052 7046 38108
rect 7046 38052 7102 38108
rect 7102 38052 7106 38108
rect 7042 38048 7106 38052
rect 7122 38108 7186 38112
rect 7122 38052 7126 38108
rect 7126 38052 7182 38108
rect 7182 38052 7186 38108
rect 7122 38048 7186 38052
rect 12813 38108 12877 38112
rect 12813 38052 12817 38108
rect 12817 38052 12873 38108
rect 12873 38052 12877 38108
rect 12813 38048 12877 38052
rect 12893 38108 12957 38112
rect 12893 38052 12897 38108
rect 12897 38052 12953 38108
rect 12953 38052 12957 38108
rect 12893 38048 12957 38052
rect 12973 38108 13037 38112
rect 12973 38052 12977 38108
rect 12977 38052 13033 38108
rect 13033 38052 13037 38108
rect 12973 38048 13037 38052
rect 13053 38108 13117 38112
rect 13053 38052 13057 38108
rect 13057 38052 13113 38108
rect 13113 38052 13117 38108
rect 13053 38048 13117 38052
rect 3917 37564 3981 37568
rect 3917 37508 3921 37564
rect 3921 37508 3977 37564
rect 3977 37508 3981 37564
rect 3917 37504 3981 37508
rect 3997 37564 4061 37568
rect 3997 37508 4001 37564
rect 4001 37508 4057 37564
rect 4057 37508 4061 37564
rect 3997 37504 4061 37508
rect 4077 37564 4141 37568
rect 4077 37508 4081 37564
rect 4081 37508 4137 37564
rect 4137 37508 4141 37564
rect 4077 37504 4141 37508
rect 4157 37564 4221 37568
rect 4157 37508 4161 37564
rect 4161 37508 4217 37564
rect 4217 37508 4221 37564
rect 4157 37504 4221 37508
rect 9848 37564 9912 37568
rect 9848 37508 9852 37564
rect 9852 37508 9908 37564
rect 9908 37508 9912 37564
rect 9848 37504 9912 37508
rect 9928 37564 9992 37568
rect 9928 37508 9932 37564
rect 9932 37508 9988 37564
rect 9988 37508 9992 37564
rect 9928 37504 9992 37508
rect 10008 37564 10072 37568
rect 10008 37508 10012 37564
rect 10012 37508 10068 37564
rect 10068 37508 10072 37564
rect 10008 37504 10072 37508
rect 10088 37564 10152 37568
rect 10088 37508 10092 37564
rect 10092 37508 10148 37564
rect 10148 37508 10152 37564
rect 10088 37504 10152 37508
rect 15778 37564 15842 37568
rect 15778 37508 15782 37564
rect 15782 37508 15838 37564
rect 15838 37508 15842 37564
rect 15778 37504 15842 37508
rect 15858 37564 15922 37568
rect 15858 37508 15862 37564
rect 15862 37508 15918 37564
rect 15918 37508 15922 37564
rect 15858 37504 15922 37508
rect 15938 37564 16002 37568
rect 15938 37508 15942 37564
rect 15942 37508 15998 37564
rect 15998 37508 16002 37564
rect 15938 37504 16002 37508
rect 16018 37564 16082 37568
rect 16018 37508 16022 37564
rect 16022 37508 16078 37564
rect 16078 37508 16082 37564
rect 16018 37504 16082 37508
rect 6882 37020 6946 37024
rect 6882 36964 6886 37020
rect 6886 36964 6942 37020
rect 6942 36964 6946 37020
rect 6882 36960 6946 36964
rect 6962 37020 7026 37024
rect 6962 36964 6966 37020
rect 6966 36964 7022 37020
rect 7022 36964 7026 37020
rect 6962 36960 7026 36964
rect 7042 37020 7106 37024
rect 7042 36964 7046 37020
rect 7046 36964 7102 37020
rect 7102 36964 7106 37020
rect 7042 36960 7106 36964
rect 7122 37020 7186 37024
rect 7122 36964 7126 37020
rect 7126 36964 7182 37020
rect 7182 36964 7186 37020
rect 7122 36960 7186 36964
rect 12813 37020 12877 37024
rect 12813 36964 12817 37020
rect 12817 36964 12873 37020
rect 12873 36964 12877 37020
rect 12813 36960 12877 36964
rect 12893 37020 12957 37024
rect 12893 36964 12897 37020
rect 12897 36964 12953 37020
rect 12953 36964 12957 37020
rect 12893 36960 12957 36964
rect 12973 37020 13037 37024
rect 12973 36964 12977 37020
rect 12977 36964 13033 37020
rect 13033 36964 13037 37020
rect 12973 36960 13037 36964
rect 13053 37020 13117 37024
rect 13053 36964 13057 37020
rect 13057 36964 13113 37020
rect 13113 36964 13117 37020
rect 13053 36960 13117 36964
rect 3917 36476 3981 36480
rect 3917 36420 3921 36476
rect 3921 36420 3977 36476
rect 3977 36420 3981 36476
rect 3917 36416 3981 36420
rect 3997 36476 4061 36480
rect 3997 36420 4001 36476
rect 4001 36420 4057 36476
rect 4057 36420 4061 36476
rect 3997 36416 4061 36420
rect 4077 36476 4141 36480
rect 4077 36420 4081 36476
rect 4081 36420 4137 36476
rect 4137 36420 4141 36476
rect 4077 36416 4141 36420
rect 4157 36476 4221 36480
rect 4157 36420 4161 36476
rect 4161 36420 4217 36476
rect 4217 36420 4221 36476
rect 4157 36416 4221 36420
rect 9848 36476 9912 36480
rect 9848 36420 9852 36476
rect 9852 36420 9908 36476
rect 9908 36420 9912 36476
rect 9848 36416 9912 36420
rect 9928 36476 9992 36480
rect 9928 36420 9932 36476
rect 9932 36420 9988 36476
rect 9988 36420 9992 36476
rect 9928 36416 9992 36420
rect 10008 36476 10072 36480
rect 10008 36420 10012 36476
rect 10012 36420 10068 36476
rect 10068 36420 10072 36476
rect 10008 36416 10072 36420
rect 10088 36476 10152 36480
rect 10088 36420 10092 36476
rect 10092 36420 10148 36476
rect 10148 36420 10152 36476
rect 10088 36416 10152 36420
rect 15778 36476 15842 36480
rect 15778 36420 15782 36476
rect 15782 36420 15838 36476
rect 15838 36420 15842 36476
rect 15778 36416 15842 36420
rect 15858 36476 15922 36480
rect 15858 36420 15862 36476
rect 15862 36420 15918 36476
rect 15918 36420 15922 36476
rect 15858 36416 15922 36420
rect 15938 36476 16002 36480
rect 15938 36420 15942 36476
rect 15942 36420 15998 36476
rect 15998 36420 16002 36476
rect 15938 36416 16002 36420
rect 16018 36476 16082 36480
rect 16018 36420 16022 36476
rect 16022 36420 16078 36476
rect 16078 36420 16082 36476
rect 16018 36416 16082 36420
rect 6882 35932 6946 35936
rect 6882 35876 6886 35932
rect 6886 35876 6942 35932
rect 6942 35876 6946 35932
rect 6882 35872 6946 35876
rect 6962 35932 7026 35936
rect 6962 35876 6966 35932
rect 6966 35876 7022 35932
rect 7022 35876 7026 35932
rect 6962 35872 7026 35876
rect 7042 35932 7106 35936
rect 7042 35876 7046 35932
rect 7046 35876 7102 35932
rect 7102 35876 7106 35932
rect 7042 35872 7106 35876
rect 7122 35932 7186 35936
rect 7122 35876 7126 35932
rect 7126 35876 7182 35932
rect 7182 35876 7186 35932
rect 7122 35872 7186 35876
rect 12813 35932 12877 35936
rect 12813 35876 12817 35932
rect 12817 35876 12873 35932
rect 12873 35876 12877 35932
rect 12813 35872 12877 35876
rect 12893 35932 12957 35936
rect 12893 35876 12897 35932
rect 12897 35876 12953 35932
rect 12953 35876 12957 35932
rect 12893 35872 12957 35876
rect 12973 35932 13037 35936
rect 12973 35876 12977 35932
rect 12977 35876 13033 35932
rect 13033 35876 13037 35932
rect 12973 35872 13037 35876
rect 13053 35932 13117 35936
rect 13053 35876 13057 35932
rect 13057 35876 13113 35932
rect 13113 35876 13117 35932
rect 13053 35872 13117 35876
rect 3917 35388 3981 35392
rect 3917 35332 3921 35388
rect 3921 35332 3977 35388
rect 3977 35332 3981 35388
rect 3917 35328 3981 35332
rect 3997 35388 4061 35392
rect 3997 35332 4001 35388
rect 4001 35332 4057 35388
rect 4057 35332 4061 35388
rect 3997 35328 4061 35332
rect 4077 35388 4141 35392
rect 4077 35332 4081 35388
rect 4081 35332 4137 35388
rect 4137 35332 4141 35388
rect 4077 35328 4141 35332
rect 4157 35388 4221 35392
rect 4157 35332 4161 35388
rect 4161 35332 4217 35388
rect 4217 35332 4221 35388
rect 4157 35328 4221 35332
rect 9848 35388 9912 35392
rect 9848 35332 9852 35388
rect 9852 35332 9908 35388
rect 9908 35332 9912 35388
rect 9848 35328 9912 35332
rect 9928 35388 9992 35392
rect 9928 35332 9932 35388
rect 9932 35332 9988 35388
rect 9988 35332 9992 35388
rect 9928 35328 9992 35332
rect 10008 35388 10072 35392
rect 10008 35332 10012 35388
rect 10012 35332 10068 35388
rect 10068 35332 10072 35388
rect 10008 35328 10072 35332
rect 10088 35388 10152 35392
rect 10088 35332 10092 35388
rect 10092 35332 10148 35388
rect 10148 35332 10152 35388
rect 10088 35328 10152 35332
rect 15778 35388 15842 35392
rect 15778 35332 15782 35388
rect 15782 35332 15838 35388
rect 15838 35332 15842 35388
rect 15778 35328 15842 35332
rect 15858 35388 15922 35392
rect 15858 35332 15862 35388
rect 15862 35332 15918 35388
rect 15918 35332 15922 35388
rect 15858 35328 15922 35332
rect 15938 35388 16002 35392
rect 15938 35332 15942 35388
rect 15942 35332 15998 35388
rect 15998 35332 16002 35388
rect 15938 35328 16002 35332
rect 16018 35388 16082 35392
rect 16018 35332 16022 35388
rect 16022 35332 16078 35388
rect 16078 35332 16082 35388
rect 16018 35328 16082 35332
rect 6882 34844 6946 34848
rect 6882 34788 6886 34844
rect 6886 34788 6942 34844
rect 6942 34788 6946 34844
rect 6882 34784 6946 34788
rect 6962 34844 7026 34848
rect 6962 34788 6966 34844
rect 6966 34788 7022 34844
rect 7022 34788 7026 34844
rect 6962 34784 7026 34788
rect 7042 34844 7106 34848
rect 7042 34788 7046 34844
rect 7046 34788 7102 34844
rect 7102 34788 7106 34844
rect 7042 34784 7106 34788
rect 7122 34844 7186 34848
rect 7122 34788 7126 34844
rect 7126 34788 7182 34844
rect 7182 34788 7186 34844
rect 7122 34784 7186 34788
rect 12813 34844 12877 34848
rect 12813 34788 12817 34844
rect 12817 34788 12873 34844
rect 12873 34788 12877 34844
rect 12813 34784 12877 34788
rect 12893 34844 12957 34848
rect 12893 34788 12897 34844
rect 12897 34788 12953 34844
rect 12953 34788 12957 34844
rect 12893 34784 12957 34788
rect 12973 34844 13037 34848
rect 12973 34788 12977 34844
rect 12977 34788 13033 34844
rect 13033 34788 13037 34844
rect 12973 34784 13037 34788
rect 13053 34844 13117 34848
rect 13053 34788 13057 34844
rect 13057 34788 13113 34844
rect 13113 34788 13117 34844
rect 13053 34784 13117 34788
rect 3917 34300 3981 34304
rect 3917 34244 3921 34300
rect 3921 34244 3977 34300
rect 3977 34244 3981 34300
rect 3917 34240 3981 34244
rect 3997 34300 4061 34304
rect 3997 34244 4001 34300
rect 4001 34244 4057 34300
rect 4057 34244 4061 34300
rect 3997 34240 4061 34244
rect 4077 34300 4141 34304
rect 4077 34244 4081 34300
rect 4081 34244 4137 34300
rect 4137 34244 4141 34300
rect 4077 34240 4141 34244
rect 4157 34300 4221 34304
rect 4157 34244 4161 34300
rect 4161 34244 4217 34300
rect 4217 34244 4221 34300
rect 4157 34240 4221 34244
rect 9848 34300 9912 34304
rect 9848 34244 9852 34300
rect 9852 34244 9908 34300
rect 9908 34244 9912 34300
rect 9848 34240 9912 34244
rect 9928 34300 9992 34304
rect 9928 34244 9932 34300
rect 9932 34244 9988 34300
rect 9988 34244 9992 34300
rect 9928 34240 9992 34244
rect 10008 34300 10072 34304
rect 10008 34244 10012 34300
rect 10012 34244 10068 34300
rect 10068 34244 10072 34300
rect 10008 34240 10072 34244
rect 10088 34300 10152 34304
rect 10088 34244 10092 34300
rect 10092 34244 10148 34300
rect 10148 34244 10152 34300
rect 10088 34240 10152 34244
rect 15778 34300 15842 34304
rect 15778 34244 15782 34300
rect 15782 34244 15838 34300
rect 15838 34244 15842 34300
rect 15778 34240 15842 34244
rect 15858 34300 15922 34304
rect 15858 34244 15862 34300
rect 15862 34244 15918 34300
rect 15918 34244 15922 34300
rect 15858 34240 15922 34244
rect 15938 34300 16002 34304
rect 15938 34244 15942 34300
rect 15942 34244 15998 34300
rect 15998 34244 16002 34300
rect 15938 34240 16002 34244
rect 16018 34300 16082 34304
rect 16018 34244 16022 34300
rect 16022 34244 16078 34300
rect 16078 34244 16082 34300
rect 16018 34240 16082 34244
rect 6882 33756 6946 33760
rect 6882 33700 6886 33756
rect 6886 33700 6942 33756
rect 6942 33700 6946 33756
rect 6882 33696 6946 33700
rect 6962 33756 7026 33760
rect 6962 33700 6966 33756
rect 6966 33700 7022 33756
rect 7022 33700 7026 33756
rect 6962 33696 7026 33700
rect 7042 33756 7106 33760
rect 7042 33700 7046 33756
rect 7046 33700 7102 33756
rect 7102 33700 7106 33756
rect 7042 33696 7106 33700
rect 7122 33756 7186 33760
rect 7122 33700 7126 33756
rect 7126 33700 7182 33756
rect 7182 33700 7186 33756
rect 7122 33696 7186 33700
rect 12813 33756 12877 33760
rect 12813 33700 12817 33756
rect 12817 33700 12873 33756
rect 12873 33700 12877 33756
rect 12813 33696 12877 33700
rect 12893 33756 12957 33760
rect 12893 33700 12897 33756
rect 12897 33700 12953 33756
rect 12953 33700 12957 33756
rect 12893 33696 12957 33700
rect 12973 33756 13037 33760
rect 12973 33700 12977 33756
rect 12977 33700 13033 33756
rect 13033 33700 13037 33756
rect 12973 33696 13037 33700
rect 13053 33756 13117 33760
rect 13053 33700 13057 33756
rect 13057 33700 13113 33756
rect 13113 33700 13117 33756
rect 13053 33696 13117 33700
rect 16620 33280 16684 33284
rect 16620 33224 16634 33280
rect 16634 33224 16684 33280
rect 16620 33220 16684 33224
rect 3917 33212 3981 33216
rect 3917 33156 3921 33212
rect 3921 33156 3977 33212
rect 3977 33156 3981 33212
rect 3917 33152 3981 33156
rect 3997 33212 4061 33216
rect 3997 33156 4001 33212
rect 4001 33156 4057 33212
rect 4057 33156 4061 33212
rect 3997 33152 4061 33156
rect 4077 33212 4141 33216
rect 4077 33156 4081 33212
rect 4081 33156 4137 33212
rect 4137 33156 4141 33212
rect 4077 33152 4141 33156
rect 4157 33212 4221 33216
rect 4157 33156 4161 33212
rect 4161 33156 4217 33212
rect 4217 33156 4221 33212
rect 4157 33152 4221 33156
rect 9848 33212 9912 33216
rect 9848 33156 9852 33212
rect 9852 33156 9908 33212
rect 9908 33156 9912 33212
rect 9848 33152 9912 33156
rect 9928 33212 9992 33216
rect 9928 33156 9932 33212
rect 9932 33156 9988 33212
rect 9988 33156 9992 33212
rect 9928 33152 9992 33156
rect 10008 33212 10072 33216
rect 10008 33156 10012 33212
rect 10012 33156 10068 33212
rect 10068 33156 10072 33212
rect 10008 33152 10072 33156
rect 10088 33212 10152 33216
rect 10088 33156 10092 33212
rect 10092 33156 10148 33212
rect 10148 33156 10152 33212
rect 10088 33152 10152 33156
rect 15778 33212 15842 33216
rect 15778 33156 15782 33212
rect 15782 33156 15838 33212
rect 15838 33156 15842 33212
rect 15778 33152 15842 33156
rect 15858 33212 15922 33216
rect 15858 33156 15862 33212
rect 15862 33156 15918 33212
rect 15918 33156 15922 33212
rect 15858 33152 15922 33156
rect 15938 33212 16002 33216
rect 15938 33156 15942 33212
rect 15942 33156 15998 33212
rect 15998 33156 16002 33212
rect 15938 33152 16002 33156
rect 16018 33212 16082 33216
rect 16018 33156 16022 33212
rect 16022 33156 16078 33212
rect 16078 33156 16082 33212
rect 16018 33152 16082 33156
rect 6882 32668 6946 32672
rect 6882 32612 6886 32668
rect 6886 32612 6942 32668
rect 6942 32612 6946 32668
rect 6882 32608 6946 32612
rect 6962 32668 7026 32672
rect 6962 32612 6966 32668
rect 6966 32612 7022 32668
rect 7022 32612 7026 32668
rect 6962 32608 7026 32612
rect 7042 32668 7106 32672
rect 7042 32612 7046 32668
rect 7046 32612 7102 32668
rect 7102 32612 7106 32668
rect 7042 32608 7106 32612
rect 7122 32668 7186 32672
rect 7122 32612 7126 32668
rect 7126 32612 7182 32668
rect 7182 32612 7186 32668
rect 7122 32608 7186 32612
rect 12813 32668 12877 32672
rect 12813 32612 12817 32668
rect 12817 32612 12873 32668
rect 12873 32612 12877 32668
rect 12813 32608 12877 32612
rect 12893 32668 12957 32672
rect 12893 32612 12897 32668
rect 12897 32612 12953 32668
rect 12953 32612 12957 32668
rect 12893 32608 12957 32612
rect 12973 32668 13037 32672
rect 12973 32612 12977 32668
rect 12977 32612 13033 32668
rect 13033 32612 13037 32668
rect 12973 32608 13037 32612
rect 13053 32668 13117 32672
rect 13053 32612 13057 32668
rect 13057 32612 13113 32668
rect 13113 32612 13117 32668
rect 13053 32608 13117 32612
rect 3917 32124 3981 32128
rect 3917 32068 3921 32124
rect 3921 32068 3977 32124
rect 3977 32068 3981 32124
rect 3917 32064 3981 32068
rect 3997 32124 4061 32128
rect 3997 32068 4001 32124
rect 4001 32068 4057 32124
rect 4057 32068 4061 32124
rect 3997 32064 4061 32068
rect 4077 32124 4141 32128
rect 4077 32068 4081 32124
rect 4081 32068 4137 32124
rect 4137 32068 4141 32124
rect 4077 32064 4141 32068
rect 4157 32124 4221 32128
rect 4157 32068 4161 32124
rect 4161 32068 4217 32124
rect 4217 32068 4221 32124
rect 4157 32064 4221 32068
rect 9848 32124 9912 32128
rect 9848 32068 9852 32124
rect 9852 32068 9908 32124
rect 9908 32068 9912 32124
rect 9848 32064 9912 32068
rect 9928 32124 9992 32128
rect 9928 32068 9932 32124
rect 9932 32068 9988 32124
rect 9988 32068 9992 32124
rect 9928 32064 9992 32068
rect 10008 32124 10072 32128
rect 10008 32068 10012 32124
rect 10012 32068 10068 32124
rect 10068 32068 10072 32124
rect 10008 32064 10072 32068
rect 10088 32124 10152 32128
rect 10088 32068 10092 32124
rect 10092 32068 10148 32124
rect 10148 32068 10152 32124
rect 10088 32064 10152 32068
rect 15778 32124 15842 32128
rect 15778 32068 15782 32124
rect 15782 32068 15838 32124
rect 15838 32068 15842 32124
rect 15778 32064 15842 32068
rect 15858 32124 15922 32128
rect 15858 32068 15862 32124
rect 15862 32068 15918 32124
rect 15918 32068 15922 32124
rect 15858 32064 15922 32068
rect 15938 32124 16002 32128
rect 15938 32068 15942 32124
rect 15942 32068 15998 32124
rect 15998 32068 16002 32124
rect 15938 32064 16002 32068
rect 16018 32124 16082 32128
rect 16018 32068 16022 32124
rect 16022 32068 16078 32124
rect 16078 32068 16082 32124
rect 16018 32064 16082 32068
rect 6882 31580 6946 31584
rect 6882 31524 6886 31580
rect 6886 31524 6942 31580
rect 6942 31524 6946 31580
rect 6882 31520 6946 31524
rect 6962 31580 7026 31584
rect 6962 31524 6966 31580
rect 6966 31524 7022 31580
rect 7022 31524 7026 31580
rect 6962 31520 7026 31524
rect 7042 31580 7106 31584
rect 7042 31524 7046 31580
rect 7046 31524 7102 31580
rect 7102 31524 7106 31580
rect 7042 31520 7106 31524
rect 7122 31580 7186 31584
rect 7122 31524 7126 31580
rect 7126 31524 7182 31580
rect 7182 31524 7186 31580
rect 7122 31520 7186 31524
rect 12813 31580 12877 31584
rect 12813 31524 12817 31580
rect 12817 31524 12873 31580
rect 12873 31524 12877 31580
rect 12813 31520 12877 31524
rect 12893 31580 12957 31584
rect 12893 31524 12897 31580
rect 12897 31524 12953 31580
rect 12953 31524 12957 31580
rect 12893 31520 12957 31524
rect 12973 31580 13037 31584
rect 12973 31524 12977 31580
rect 12977 31524 13033 31580
rect 13033 31524 13037 31580
rect 12973 31520 13037 31524
rect 13053 31580 13117 31584
rect 13053 31524 13057 31580
rect 13057 31524 13113 31580
rect 13113 31524 13117 31580
rect 13053 31520 13117 31524
rect 3917 31036 3981 31040
rect 3917 30980 3921 31036
rect 3921 30980 3977 31036
rect 3977 30980 3981 31036
rect 3917 30976 3981 30980
rect 3997 31036 4061 31040
rect 3997 30980 4001 31036
rect 4001 30980 4057 31036
rect 4057 30980 4061 31036
rect 3997 30976 4061 30980
rect 4077 31036 4141 31040
rect 4077 30980 4081 31036
rect 4081 30980 4137 31036
rect 4137 30980 4141 31036
rect 4077 30976 4141 30980
rect 4157 31036 4221 31040
rect 4157 30980 4161 31036
rect 4161 30980 4217 31036
rect 4217 30980 4221 31036
rect 4157 30976 4221 30980
rect 9848 31036 9912 31040
rect 9848 30980 9852 31036
rect 9852 30980 9908 31036
rect 9908 30980 9912 31036
rect 9848 30976 9912 30980
rect 9928 31036 9992 31040
rect 9928 30980 9932 31036
rect 9932 30980 9988 31036
rect 9988 30980 9992 31036
rect 9928 30976 9992 30980
rect 10008 31036 10072 31040
rect 10008 30980 10012 31036
rect 10012 30980 10068 31036
rect 10068 30980 10072 31036
rect 10008 30976 10072 30980
rect 10088 31036 10152 31040
rect 10088 30980 10092 31036
rect 10092 30980 10148 31036
rect 10148 30980 10152 31036
rect 10088 30976 10152 30980
rect 15778 31036 15842 31040
rect 15778 30980 15782 31036
rect 15782 30980 15838 31036
rect 15838 30980 15842 31036
rect 15778 30976 15842 30980
rect 15858 31036 15922 31040
rect 15858 30980 15862 31036
rect 15862 30980 15918 31036
rect 15918 30980 15922 31036
rect 15858 30976 15922 30980
rect 15938 31036 16002 31040
rect 15938 30980 15942 31036
rect 15942 30980 15998 31036
rect 15998 30980 16002 31036
rect 15938 30976 16002 30980
rect 16018 31036 16082 31040
rect 16018 30980 16022 31036
rect 16022 30980 16078 31036
rect 16078 30980 16082 31036
rect 16018 30976 16082 30980
rect 6882 30492 6946 30496
rect 6882 30436 6886 30492
rect 6886 30436 6942 30492
rect 6942 30436 6946 30492
rect 6882 30432 6946 30436
rect 6962 30492 7026 30496
rect 6962 30436 6966 30492
rect 6966 30436 7022 30492
rect 7022 30436 7026 30492
rect 6962 30432 7026 30436
rect 7042 30492 7106 30496
rect 7042 30436 7046 30492
rect 7046 30436 7102 30492
rect 7102 30436 7106 30492
rect 7042 30432 7106 30436
rect 7122 30492 7186 30496
rect 7122 30436 7126 30492
rect 7126 30436 7182 30492
rect 7182 30436 7186 30492
rect 7122 30432 7186 30436
rect 12813 30492 12877 30496
rect 12813 30436 12817 30492
rect 12817 30436 12873 30492
rect 12873 30436 12877 30492
rect 12813 30432 12877 30436
rect 12893 30492 12957 30496
rect 12893 30436 12897 30492
rect 12897 30436 12953 30492
rect 12953 30436 12957 30492
rect 12893 30432 12957 30436
rect 12973 30492 13037 30496
rect 12973 30436 12977 30492
rect 12977 30436 13033 30492
rect 13033 30436 13037 30492
rect 12973 30432 13037 30436
rect 13053 30492 13117 30496
rect 13053 30436 13057 30492
rect 13057 30436 13113 30492
rect 13113 30436 13117 30492
rect 13053 30432 13117 30436
rect 3917 29948 3981 29952
rect 3917 29892 3921 29948
rect 3921 29892 3977 29948
rect 3977 29892 3981 29948
rect 3917 29888 3981 29892
rect 3997 29948 4061 29952
rect 3997 29892 4001 29948
rect 4001 29892 4057 29948
rect 4057 29892 4061 29948
rect 3997 29888 4061 29892
rect 4077 29948 4141 29952
rect 4077 29892 4081 29948
rect 4081 29892 4137 29948
rect 4137 29892 4141 29948
rect 4077 29888 4141 29892
rect 4157 29948 4221 29952
rect 4157 29892 4161 29948
rect 4161 29892 4217 29948
rect 4217 29892 4221 29948
rect 4157 29888 4221 29892
rect 9848 29948 9912 29952
rect 9848 29892 9852 29948
rect 9852 29892 9908 29948
rect 9908 29892 9912 29948
rect 9848 29888 9912 29892
rect 9928 29948 9992 29952
rect 9928 29892 9932 29948
rect 9932 29892 9988 29948
rect 9988 29892 9992 29948
rect 9928 29888 9992 29892
rect 10008 29948 10072 29952
rect 10008 29892 10012 29948
rect 10012 29892 10068 29948
rect 10068 29892 10072 29948
rect 10008 29888 10072 29892
rect 10088 29948 10152 29952
rect 10088 29892 10092 29948
rect 10092 29892 10148 29948
rect 10148 29892 10152 29948
rect 10088 29888 10152 29892
rect 15778 29948 15842 29952
rect 15778 29892 15782 29948
rect 15782 29892 15838 29948
rect 15838 29892 15842 29948
rect 15778 29888 15842 29892
rect 15858 29948 15922 29952
rect 15858 29892 15862 29948
rect 15862 29892 15918 29948
rect 15918 29892 15922 29948
rect 15858 29888 15922 29892
rect 15938 29948 16002 29952
rect 15938 29892 15942 29948
rect 15942 29892 15998 29948
rect 15998 29892 16002 29948
rect 15938 29888 16002 29892
rect 16018 29948 16082 29952
rect 16018 29892 16022 29948
rect 16022 29892 16078 29948
rect 16078 29892 16082 29948
rect 16018 29888 16082 29892
rect 6882 29404 6946 29408
rect 6882 29348 6886 29404
rect 6886 29348 6942 29404
rect 6942 29348 6946 29404
rect 6882 29344 6946 29348
rect 6962 29404 7026 29408
rect 6962 29348 6966 29404
rect 6966 29348 7022 29404
rect 7022 29348 7026 29404
rect 6962 29344 7026 29348
rect 7042 29404 7106 29408
rect 7042 29348 7046 29404
rect 7046 29348 7102 29404
rect 7102 29348 7106 29404
rect 7042 29344 7106 29348
rect 7122 29404 7186 29408
rect 7122 29348 7126 29404
rect 7126 29348 7182 29404
rect 7182 29348 7186 29404
rect 7122 29344 7186 29348
rect 12813 29404 12877 29408
rect 12813 29348 12817 29404
rect 12817 29348 12873 29404
rect 12873 29348 12877 29404
rect 12813 29344 12877 29348
rect 12893 29404 12957 29408
rect 12893 29348 12897 29404
rect 12897 29348 12953 29404
rect 12953 29348 12957 29404
rect 12893 29344 12957 29348
rect 12973 29404 13037 29408
rect 12973 29348 12977 29404
rect 12977 29348 13033 29404
rect 13033 29348 13037 29404
rect 12973 29344 13037 29348
rect 13053 29404 13117 29408
rect 13053 29348 13057 29404
rect 13057 29348 13113 29404
rect 13113 29348 13117 29404
rect 13053 29344 13117 29348
rect 3917 28860 3981 28864
rect 3917 28804 3921 28860
rect 3921 28804 3977 28860
rect 3977 28804 3981 28860
rect 3917 28800 3981 28804
rect 3997 28860 4061 28864
rect 3997 28804 4001 28860
rect 4001 28804 4057 28860
rect 4057 28804 4061 28860
rect 3997 28800 4061 28804
rect 4077 28860 4141 28864
rect 4077 28804 4081 28860
rect 4081 28804 4137 28860
rect 4137 28804 4141 28860
rect 4077 28800 4141 28804
rect 4157 28860 4221 28864
rect 4157 28804 4161 28860
rect 4161 28804 4217 28860
rect 4217 28804 4221 28860
rect 4157 28800 4221 28804
rect 9848 28860 9912 28864
rect 9848 28804 9852 28860
rect 9852 28804 9908 28860
rect 9908 28804 9912 28860
rect 9848 28800 9912 28804
rect 9928 28860 9992 28864
rect 9928 28804 9932 28860
rect 9932 28804 9988 28860
rect 9988 28804 9992 28860
rect 9928 28800 9992 28804
rect 10008 28860 10072 28864
rect 10008 28804 10012 28860
rect 10012 28804 10068 28860
rect 10068 28804 10072 28860
rect 10008 28800 10072 28804
rect 10088 28860 10152 28864
rect 10088 28804 10092 28860
rect 10092 28804 10148 28860
rect 10148 28804 10152 28860
rect 10088 28800 10152 28804
rect 15778 28860 15842 28864
rect 15778 28804 15782 28860
rect 15782 28804 15838 28860
rect 15838 28804 15842 28860
rect 15778 28800 15842 28804
rect 15858 28860 15922 28864
rect 15858 28804 15862 28860
rect 15862 28804 15918 28860
rect 15918 28804 15922 28860
rect 15858 28800 15922 28804
rect 15938 28860 16002 28864
rect 15938 28804 15942 28860
rect 15942 28804 15998 28860
rect 15998 28804 16002 28860
rect 15938 28800 16002 28804
rect 16018 28860 16082 28864
rect 16018 28804 16022 28860
rect 16022 28804 16078 28860
rect 16078 28804 16082 28860
rect 16018 28800 16082 28804
rect 6882 28316 6946 28320
rect 6882 28260 6886 28316
rect 6886 28260 6942 28316
rect 6942 28260 6946 28316
rect 6882 28256 6946 28260
rect 6962 28316 7026 28320
rect 6962 28260 6966 28316
rect 6966 28260 7022 28316
rect 7022 28260 7026 28316
rect 6962 28256 7026 28260
rect 7042 28316 7106 28320
rect 7042 28260 7046 28316
rect 7046 28260 7102 28316
rect 7102 28260 7106 28316
rect 7042 28256 7106 28260
rect 7122 28316 7186 28320
rect 7122 28260 7126 28316
rect 7126 28260 7182 28316
rect 7182 28260 7186 28316
rect 7122 28256 7186 28260
rect 12813 28316 12877 28320
rect 12813 28260 12817 28316
rect 12817 28260 12873 28316
rect 12873 28260 12877 28316
rect 12813 28256 12877 28260
rect 12893 28316 12957 28320
rect 12893 28260 12897 28316
rect 12897 28260 12953 28316
rect 12953 28260 12957 28316
rect 12893 28256 12957 28260
rect 12973 28316 13037 28320
rect 12973 28260 12977 28316
rect 12977 28260 13033 28316
rect 13033 28260 13037 28316
rect 12973 28256 13037 28260
rect 13053 28316 13117 28320
rect 13053 28260 13057 28316
rect 13057 28260 13113 28316
rect 13113 28260 13117 28316
rect 13053 28256 13117 28260
rect 3917 27772 3981 27776
rect 3917 27716 3921 27772
rect 3921 27716 3977 27772
rect 3977 27716 3981 27772
rect 3917 27712 3981 27716
rect 3997 27772 4061 27776
rect 3997 27716 4001 27772
rect 4001 27716 4057 27772
rect 4057 27716 4061 27772
rect 3997 27712 4061 27716
rect 4077 27772 4141 27776
rect 4077 27716 4081 27772
rect 4081 27716 4137 27772
rect 4137 27716 4141 27772
rect 4077 27712 4141 27716
rect 4157 27772 4221 27776
rect 4157 27716 4161 27772
rect 4161 27716 4217 27772
rect 4217 27716 4221 27772
rect 4157 27712 4221 27716
rect 9848 27772 9912 27776
rect 9848 27716 9852 27772
rect 9852 27716 9908 27772
rect 9908 27716 9912 27772
rect 9848 27712 9912 27716
rect 9928 27772 9992 27776
rect 9928 27716 9932 27772
rect 9932 27716 9988 27772
rect 9988 27716 9992 27772
rect 9928 27712 9992 27716
rect 10008 27772 10072 27776
rect 10008 27716 10012 27772
rect 10012 27716 10068 27772
rect 10068 27716 10072 27772
rect 10008 27712 10072 27716
rect 10088 27772 10152 27776
rect 10088 27716 10092 27772
rect 10092 27716 10148 27772
rect 10148 27716 10152 27772
rect 10088 27712 10152 27716
rect 15778 27772 15842 27776
rect 15778 27716 15782 27772
rect 15782 27716 15838 27772
rect 15838 27716 15842 27772
rect 15778 27712 15842 27716
rect 15858 27772 15922 27776
rect 15858 27716 15862 27772
rect 15862 27716 15918 27772
rect 15918 27716 15922 27772
rect 15858 27712 15922 27716
rect 15938 27772 16002 27776
rect 15938 27716 15942 27772
rect 15942 27716 15998 27772
rect 15998 27716 16002 27772
rect 15938 27712 16002 27716
rect 16018 27772 16082 27776
rect 16018 27716 16022 27772
rect 16022 27716 16078 27772
rect 16078 27716 16082 27772
rect 16018 27712 16082 27716
rect 6882 27228 6946 27232
rect 6882 27172 6886 27228
rect 6886 27172 6942 27228
rect 6942 27172 6946 27228
rect 6882 27168 6946 27172
rect 6962 27228 7026 27232
rect 6962 27172 6966 27228
rect 6966 27172 7022 27228
rect 7022 27172 7026 27228
rect 6962 27168 7026 27172
rect 7042 27228 7106 27232
rect 7042 27172 7046 27228
rect 7046 27172 7102 27228
rect 7102 27172 7106 27228
rect 7042 27168 7106 27172
rect 7122 27228 7186 27232
rect 7122 27172 7126 27228
rect 7126 27172 7182 27228
rect 7182 27172 7186 27228
rect 7122 27168 7186 27172
rect 12813 27228 12877 27232
rect 12813 27172 12817 27228
rect 12817 27172 12873 27228
rect 12873 27172 12877 27228
rect 12813 27168 12877 27172
rect 12893 27228 12957 27232
rect 12893 27172 12897 27228
rect 12897 27172 12953 27228
rect 12953 27172 12957 27228
rect 12893 27168 12957 27172
rect 12973 27228 13037 27232
rect 12973 27172 12977 27228
rect 12977 27172 13033 27228
rect 13033 27172 13037 27228
rect 12973 27168 13037 27172
rect 13053 27228 13117 27232
rect 13053 27172 13057 27228
rect 13057 27172 13113 27228
rect 13113 27172 13117 27228
rect 13053 27168 13117 27172
rect 3917 26684 3981 26688
rect 3917 26628 3921 26684
rect 3921 26628 3977 26684
rect 3977 26628 3981 26684
rect 3917 26624 3981 26628
rect 3997 26684 4061 26688
rect 3997 26628 4001 26684
rect 4001 26628 4057 26684
rect 4057 26628 4061 26684
rect 3997 26624 4061 26628
rect 4077 26684 4141 26688
rect 4077 26628 4081 26684
rect 4081 26628 4137 26684
rect 4137 26628 4141 26684
rect 4077 26624 4141 26628
rect 4157 26684 4221 26688
rect 4157 26628 4161 26684
rect 4161 26628 4217 26684
rect 4217 26628 4221 26684
rect 4157 26624 4221 26628
rect 9848 26684 9912 26688
rect 9848 26628 9852 26684
rect 9852 26628 9908 26684
rect 9908 26628 9912 26684
rect 9848 26624 9912 26628
rect 9928 26684 9992 26688
rect 9928 26628 9932 26684
rect 9932 26628 9988 26684
rect 9988 26628 9992 26684
rect 9928 26624 9992 26628
rect 10008 26684 10072 26688
rect 10008 26628 10012 26684
rect 10012 26628 10068 26684
rect 10068 26628 10072 26684
rect 10008 26624 10072 26628
rect 10088 26684 10152 26688
rect 10088 26628 10092 26684
rect 10092 26628 10148 26684
rect 10148 26628 10152 26684
rect 10088 26624 10152 26628
rect 15778 26684 15842 26688
rect 15778 26628 15782 26684
rect 15782 26628 15838 26684
rect 15838 26628 15842 26684
rect 15778 26624 15842 26628
rect 15858 26684 15922 26688
rect 15858 26628 15862 26684
rect 15862 26628 15918 26684
rect 15918 26628 15922 26684
rect 15858 26624 15922 26628
rect 15938 26684 16002 26688
rect 15938 26628 15942 26684
rect 15942 26628 15998 26684
rect 15998 26628 16002 26684
rect 15938 26624 16002 26628
rect 16018 26684 16082 26688
rect 16018 26628 16022 26684
rect 16022 26628 16078 26684
rect 16078 26628 16082 26684
rect 16018 26624 16082 26628
rect 6882 26140 6946 26144
rect 6882 26084 6886 26140
rect 6886 26084 6942 26140
rect 6942 26084 6946 26140
rect 6882 26080 6946 26084
rect 6962 26140 7026 26144
rect 6962 26084 6966 26140
rect 6966 26084 7022 26140
rect 7022 26084 7026 26140
rect 6962 26080 7026 26084
rect 7042 26140 7106 26144
rect 7042 26084 7046 26140
rect 7046 26084 7102 26140
rect 7102 26084 7106 26140
rect 7042 26080 7106 26084
rect 7122 26140 7186 26144
rect 7122 26084 7126 26140
rect 7126 26084 7182 26140
rect 7182 26084 7186 26140
rect 7122 26080 7186 26084
rect 12813 26140 12877 26144
rect 12813 26084 12817 26140
rect 12817 26084 12873 26140
rect 12873 26084 12877 26140
rect 12813 26080 12877 26084
rect 12893 26140 12957 26144
rect 12893 26084 12897 26140
rect 12897 26084 12953 26140
rect 12953 26084 12957 26140
rect 12893 26080 12957 26084
rect 12973 26140 13037 26144
rect 12973 26084 12977 26140
rect 12977 26084 13033 26140
rect 13033 26084 13037 26140
rect 12973 26080 13037 26084
rect 13053 26140 13117 26144
rect 13053 26084 13057 26140
rect 13057 26084 13113 26140
rect 13113 26084 13117 26140
rect 13053 26080 13117 26084
rect 3917 25596 3981 25600
rect 3917 25540 3921 25596
rect 3921 25540 3977 25596
rect 3977 25540 3981 25596
rect 3917 25536 3981 25540
rect 3997 25596 4061 25600
rect 3997 25540 4001 25596
rect 4001 25540 4057 25596
rect 4057 25540 4061 25596
rect 3997 25536 4061 25540
rect 4077 25596 4141 25600
rect 4077 25540 4081 25596
rect 4081 25540 4137 25596
rect 4137 25540 4141 25596
rect 4077 25536 4141 25540
rect 4157 25596 4221 25600
rect 4157 25540 4161 25596
rect 4161 25540 4217 25596
rect 4217 25540 4221 25596
rect 4157 25536 4221 25540
rect 9848 25596 9912 25600
rect 9848 25540 9852 25596
rect 9852 25540 9908 25596
rect 9908 25540 9912 25596
rect 9848 25536 9912 25540
rect 9928 25596 9992 25600
rect 9928 25540 9932 25596
rect 9932 25540 9988 25596
rect 9988 25540 9992 25596
rect 9928 25536 9992 25540
rect 10008 25596 10072 25600
rect 10008 25540 10012 25596
rect 10012 25540 10068 25596
rect 10068 25540 10072 25596
rect 10008 25536 10072 25540
rect 10088 25596 10152 25600
rect 10088 25540 10092 25596
rect 10092 25540 10148 25596
rect 10148 25540 10152 25596
rect 10088 25536 10152 25540
rect 15778 25596 15842 25600
rect 15778 25540 15782 25596
rect 15782 25540 15838 25596
rect 15838 25540 15842 25596
rect 15778 25536 15842 25540
rect 15858 25596 15922 25600
rect 15858 25540 15862 25596
rect 15862 25540 15918 25596
rect 15918 25540 15922 25596
rect 15858 25536 15922 25540
rect 15938 25596 16002 25600
rect 15938 25540 15942 25596
rect 15942 25540 15998 25596
rect 15998 25540 16002 25596
rect 15938 25536 16002 25540
rect 16018 25596 16082 25600
rect 16018 25540 16022 25596
rect 16022 25540 16078 25596
rect 16078 25540 16082 25596
rect 16018 25536 16082 25540
rect 15516 25468 15580 25532
rect 6882 25052 6946 25056
rect 6882 24996 6886 25052
rect 6886 24996 6942 25052
rect 6942 24996 6946 25052
rect 6882 24992 6946 24996
rect 6962 25052 7026 25056
rect 6962 24996 6966 25052
rect 6966 24996 7022 25052
rect 7022 24996 7026 25052
rect 6962 24992 7026 24996
rect 7042 25052 7106 25056
rect 7042 24996 7046 25052
rect 7046 24996 7102 25052
rect 7102 24996 7106 25052
rect 7042 24992 7106 24996
rect 7122 25052 7186 25056
rect 7122 24996 7126 25052
rect 7126 24996 7182 25052
rect 7182 24996 7186 25052
rect 7122 24992 7186 24996
rect 12813 25052 12877 25056
rect 12813 24996 12817 25052
rect 12817 24996 12873 25052
rect 12873 24996 12877 25052
rect 12813 24992 12877 24996
rect 12893 25052 12957 25056
rect 12893 24996 12897 25052
rect 12897 24996 12953 25052
rect 12953 24996 12957 25052
rect 12893 24992 12957 24996
rect 12973 25052 13037 25056
rect 12973 24996 12977 25052
rect 12977 24996 13033 25052
rect 13033 24996 13037 25052
rect 12973 24992 13037 24996
rect 13053 25052 13117 25056
rect 13053 24996 13057 25052
rect 13057 24996 13113 25052
rect 13113 24996 13117 25052
rect 13053 24992 13117 24996
rect 3917 24508 3981 24512
rect 3917 24452 3921 24508
rect 3921 24452 3977 24508
rect 3977 24452 3981 24508
rect 3917 24448 3981 24452
rect 3997 24508 4061 24512
rect 3997 24452 4001 24508
rect 4001 24452 4057 24508
rect 4057 24452 4061 24508
rect 3997 24448 4061 24452
rect 4077 24508 4141 24512
rect 4077 24452 4081 24508
rect 4081 24452 4137 24508
rect 4137 24452 4141 24508
rect 4077 24448 4141 24452
rect 4157 24508 4221 24512
rect 4157 24452 4161 24508
rect 4161 24452 4217 24508
rect 4217 24452 4221 24508
rect 4157 24448 4221 24452
rect 9848 24508 9912 24512
rect 9848 24452 9852 24508
rect 9852 24452 9908 24508
rect 9908 24452 9912 24508
rect 9848 24448 9912 24452
rect 9928 24508 9992 24512
rect 9928 24452 9932 24508
rect 9932 24452 9988 24508
rect 9988 24452 9992 24508
rect 9928 24448 9992 24452
rect 10008 24508 10072 24512
rect 10008 24452 10012 24508
rect 10012 24452 10068 24508
rect 10068 24452 10072 24508
rect 10008 24448 10072 24452
rect 10088 24508 10152 24512
rect 10088 24452 10092 24508
rect 10092 24452 10148 24508
rect 10148 24452 10152 24508
rect 10088 24448 10152 24452
rect 15778 24508 15842 24512
rect 15778 24452 15782 24508
rect 15782 24452 15838 24508
rect 15838 24452 15842 24508
rect 15778 24448 15842 24452
rect 15858 24508 15922 24512
rect 15858 24452 15862 24508
rect 15862 24452 15918 24508
rect 15918 24452 15922 24508
rect 15858 24448 15922 24452
rect 15938 24508 16002 24512
rect 15938 24452 15942 24508
rect 15942 24452 15998 24508
rect 15998 24452 16002 24508
rect 15938 24448 16002 24452
rect 16018 24508 16082 24512
rect 16018 24452 16022 24508
rect 16022 24452 16078 24508
rect 16078 24452 16082 24508
rect 16018 24448 16082 24452
rect 6882 23964 6946 23968
rect 6882 23908 6886 23964
rect 6886 23908 6942 23964
rect 6942 23908 6946 23964
rect 6882 23904 6946 23908
rect 6962 23964 7026 23968
rect 6962 23908 6966 23964
rect 6966 23908 7022 23964
rect 7022 23908 7026 23964
rect 6962 23904 7026 23908
rect 7042 23964 7106 23968
rect 7042 23908 7046 23964
rect 7046 23908 7102 23964
rect 7102 23908 7106 23964
rect 7042 23904 7106 23908
rect 7122 23964 7186 23968
rect 7122 23908 7126 23964
rect 7126 23908 7182 23964
rect 7182 23908 7186 23964
rect 7122 23904 7186 23908
rect 12813 23964 12877 23968
rect 12813 23908 12817 23964
rect 12817 23908 12873 23964
rect 12873 23908 12877 23964
rect 12813 23904 12877 23908
rect 12893 23964 12957 23968
rect 12893 23908 12897 23964
rect 12897 23908 12953 23964
rect 12953 23908 12957 23964
rect 12893 23904 12957 23908
rect 12973 23964 13037 23968
rect 12973 23908 12977 23964
rect 12977 23908 13033 23964
rect 13033 23908 13037 23964
rect 12973 23904 13037 23908
rect 13053 23964 13117 23968
rect 13053 23908 13057 23964
rect 13057 23908 13113 23964
rect 13113 23908 13117 23964
rect 13053 23904 13117 23908
rect 3917 23420 3981 23424
rect 3917 23364 3921 23420
rect 3921 23364 3977 23420
rect 3977 23364 3981 23420
rect 3917 23360 3981 23364
rect 3997 23420 4061 23424
rect 3997 23364 4001 23420
rect 4001 23364 4057 23420
rect 4057 23364 4061 23420
rect 3997 23360 4061 23364
rect 4077 23420 4141 23424
rect 4077 23364 4081 23420
rect 4081 23364 4137 23420
rect 4137 23364 4141 23420
rect 4077 23360 4141 23364
rect 4157 23420 4221 23424
rect 4157 23364 4161 23420
rect 4161 23364 4217 23420
rect 4217 23364 4221 23420
rect 4157 23360 4221 23364
rect 9848 23420 9912 23424
rect 9848 23364 9852 23420
rect 9852 23364 9908 23420
rect 9908 23364 9912 23420
rect 9848 23360 9912 23364
rect 9928 23420 9992 23424
rect 9928 23364 9932 23420
rect 9932 23364 9988 23420
rect 9988 23364 9992 23420
rect 9928 23360 9992 23364
rect 10008 23420 10072 23424
rect 10008 23364 10012 23420
rect 10012 23364 10068 23420
rect 10068 23364 10072 23420
rect 10008 23360 10072 23364
rect 10088 23420 10152 23424
rect 10088 23364 10092 23420
rect 10092 23364 10148 23420
rect 10148 23364 10152 23420
rect 10088 23360 10152 23364
rect 15778 23420 15842 23424
rect 15778 23364 15782 23420
rect 15782 23364 15838 23420
rect 15838 23364 15842 23420
rect 15778 23360 15842 23364
rect 15858 23420 15922 23424
rect 15858 23364 15862 23420
rect 15862 23364 15918 23420
rect 15918 23364 15922 23420
rect 15858 23360 15922 23364
rect 15938 23420 16002 23424
rect 15938 23364 15942 23420
rect 15942 23364 15998 23420
rect 15998 23364 16002 23420
rect 15938 23360 16002 23364
rect 16018 23420 16082 23424
rect 16018 23364 16022 23420
rect 16022 23364 16078 23420
rect 16078 23364 16082 23420
rect 16018 23360 16082 23364
rect 6882 22876 6946 22880
rect 6882 22820 6886 22876
rect 6886 22820 6942 22876
rect 6942 22820 6946 22876
rect 6882 22816 6946 22820
rect 6962 22876 7026 22880
rect 6962 22820 6966 22876
rect 6966 22820 7022 22876
rect 7022 22820 7026 22876
rect 6962 22816 7026 22820
rect 7042 22876 7106 22880
rect 7042 22820 7046 22876
rect 7046 22820 7102 22876
rect 7102 22820 7106 22876
rect 7042 22816 7106 22820
rect 7122 22876 7186 22880
rect 7122 22820 7126 22876
rect 7126 22820 7182 22876
rect 7182 22820 7186 22876
rect 7122 22816 7186 22820
rect 12813 22876 12877 22880
rect 12813 22820 12817 22876
rect 12817 22820 12873 22876
rect 12873 22820 12877 22876
rect 12813 22816 12877 22820
rect 12893 22876 12957 22880
rect 12893 22820 12897 22876
rect 12897 22820 12953 22876
rect 12953 22820 12957 22876
rect 12893 22816 12957 22820
rect 12973 22876 13037 22880
rect 12973 22820 12977 22876
rect 12977 22820 13033 22876
rect 13033 22820 13037 22876
rect 12973 22816 13037 22820
rect 13053 22876 13117 22880
rect 13053 22820 13057 22876
rect 13057 22820 13113 22876
rect 13113 22820 13117 22876
rect 13053 22816 13117 22820
rect 3917 22332 3981 22336
rect 3917 22276 3921 22332
rect 3921 22276 3977 22332
rect 3977 22276 3981 22332
rect 3917 22272 3981 22276
rect 3997 22332 4061 22336
rect 3997 22276 4001 22332
rect 4001 22276 4057 22332
rect 4057 22276 4061 22332
rect 3997 22272 4061 22276
rect 4077 22332 4141 22336
rect 4077 22276 4081 22332
rect 4081 22276 4137 22332
rect 4137 22276 4141 22332
rect 4077 22272 4141 22276
rect 4157 22332 4221 22336
rect 4157 22276 4161 22332
rect 4161 22276 4217 22332
rect 4217 22276 4221 22332
rect 4157 22272 4221 22276
rect 9848 22332 9912 22336
rect 9848 22276 9852 22332
rect 9852 22276 9908 22332
rect 9908 22276 9912 22332
rect 9848 22272 9912 22276
rect 9928 22332 9992 22336
rect 9928 22276 9932 22332
rect 9932 22276 9988 22332
rect 9988 22276 9992 22332
rect 9928 22272 9992 22276
rect 10008 22332 10072 22336
rect 10008 22276 10012 22332
rect 10012 22276 10068 22332
rect 10068 22276 10072 22332
rect 10008 22272 10072 22276
rect 10088 22332 10152 22336
rect 10088 22276 10092 22332
rect 10092 22276 10148 22332
rect 10148 22276 10152 22332
rect 10088 22272 10152 22276
rect 15778 22332 15842 22336
rect 15778 22276 15782 22332
rect 15782 22276 15838 22332
rect 15838 22276 15842 22332
rect 15778 22272 15842 22276
rect 15858 22332 15922 22336
rect 15858 22276 15862 22332
rect 15862 22276 15918 22332
rect 15918 22276 15922 22332
rect 15858 22272 15922 22276
rect 15938 22332 16002 22336
rect 15938 22276 15942 22332
rect 15942 22276 15998 22332
rect 15998 22276 16002 22332
rect 15938 22272 16002 22276
rect 16018 22332 16082 22336
rect 16018 22276 16022 22332
rect 16022 22276 16078 22332
rect 16078 22276 16082 22332
rect 16018 22272 16082 22276
rect 6882 21788 6946 21792
rect 6882 21732 6886 21788
rect 6886 21732 6942 21788
rect 6942 21732 6946 21788
rect 6882 21728 6946 21732
rect 6962 21788 7026 21792
rect 6962 21732 6966 21788
rect 6966 21732 7022 21788
rect 7022 21732 7026 21788
rect 6962 21728 7026 21732
rect 7042 21788 7106 21792
rect 7042 21732 7046 21788
rect 7046 21732 7102 21788
rect 7102 21732 7106 21788
rect 7042 21728 7106 21732
rect 7122 21788 7186 21792
rect 7122 21732 7126 21788
rect 7126 21732 7182 21788
rect 7182 21732 7186 21788
rect 7122 21728 7186 21732
rect 12813 21788 12877 21792
rect 12813 21732 12817 21788
rect 12817 21732 12873 21788
rect 12873 21732 12877 21788
rect 12813 21728 12877 21732
rect 12893 21788 12957 21792
rect 12893 21732 12897 21788
rect 12897 21732 12953 21788
rect 12953 21732 12957 21788
rect 12893 21728 12957 21732
rect 12973 21788 13037 21792
rect 12973 21732 12977 21788
rect 12977 21732 13033 21788
rect 13033 21732 13037 21788
rect 12973 21728 13037 21732
rect 13053 21788 13117 21792
rect 13053 21732 13057 21788
rect 13057 21732 13113 21788
rect 13113 21732 13117 21788
rect 13053 21728 13117 21732
rect 3917 21244 3981 21248
rect 3917 21188 3921 21244
rect 3921 21188 3977 21244
rect 3977 21188 3981 21244
rect 3917 21184 3981 21188
rect 3997 21244 4061 21248
rect 3997 21188 4001 21244
rect 4001 21188 4057 21244
rect 4057 21188 4061 21244
rect 3997 21184 4061 21188
rect 4077 21244 4141 21248
rect 4077 21188 4081 21244
rect 4081 21188 4137 21244
rect 4137 21188 4141 21244
rect 4077 21184 4141 21188
rect 4157 21244 4221 21248
rect 4157 21188 4161 21244
rect 4161 21188 4217 21244
rect 4217 21188 4221 21244
rect 4157 21184 4221 21188
rect 9848 21244 9912 21248
rect 9848 21188 9852 21244
rect 9852 21188 9908 21244
rect 9908 21188 9912 21244
rect 9848 21184 9912 21188
rect 9928 21244 9992 21248
rect 9928 21188 9932 21244
rect 9932 21188 9988 21244
rect 9988 21188 9992 21244
rect 9928 21184 9992 21188
rect 10008 21244 10072 21248
rect 10008 21188 10012 21244
rect 10012 21188 10068 21244
rect 10068 21188 10072 21244
rect 10008 21184 10072 21188
rect 10088 21244 10152 21248
rect 10088 21188 10092 21244
rect 10092 21188 10148 21244
rect 10148 21188 10152 21244
rect 10088 21184 10152 21188
rect 15778 21244 15842 21248
rect 15778 21188 15782 21244
rect 15782 21188 15838 21244
rect 15838 21188 15842 21244
rect 15778 21184 15842 21188
rect 15858 21244 15922 21248
rect 15858 21188 15862 21244
rect 15862 21188 15918 21244
rect 15918 21188 15922 21244
rect 15858 21184 15922 21188
rect 15938 21244 16002 21248
rect 15938 21188 15942 21244
rect 15942 21188 15998 21244
rect 15998 21188 16002 21244
rect 15938 21184 16002 21188
rect 16018 21244 16082 21248
rect 16018 21188 16022 21244
rect 16022 21188 16078 21244
rect 16078 21188 16082 21244
rect 16018 21184 16082 21188
rect 6882 20700 6946 20704
rect 6882 20644 6886 20700
rect 6886 20644 6942 20700
rect 6942 20644 6946 20700
rect 6882 20640 6946 20644
rect 6962 20700 7026 20704
rect 6962 20644 6966 20700
rect 6966 20644 7022 20700
rect 7022 20644 7026 20700
rect 6962 20640 7026 20644
rect 7042 20700 7106 20704
rect 7042 20644 7046 20700
rect 7046 20644 7102 20700
rect 7102 20644 7106 20700
rect 7042 20640 7106 20644
rect 7122 20700 7186 20704
rect 7122 20644 7126 20700
rect 7126 20644 7182 20700
rect 7182 20644 7186 20700
rect 7122 20640 7186 20644
rect 12813 20700 12877 20704
rect 12813 20644 12817 20700
rect 12817 20644 12873 20700
rect 12873 20644 12877 20700
rect 12813 20640 12877 20644
rect 12893 20700 12957 20704
rect 12893 20644 12897 20700
rect 12897 20644 12953 20700
rect 12953 20644 12957 20700
rect 12893 20640 12957 20644
rect 12973 20700 13037 20704
rect 12973 20644 12977 20700
rect 12977 20644 13033 20700
rect 13033 20644 13037 20700
rect 12973 20640 13037 20644
rect 13053 20700 13117 20704
rect 13053 20644 13057 20700
rect 13057 20644 13113 20700
rect 13113 20644 13117 20700
rect 13053 20640 13117 20644
rect 3917 20156 3981 20160
rect 3917 20100 3921 20156
rect 3921 20100 3977 20156
rect 3977 20100 3981 20156
rect 3917 20096 3981 20100
rect 3997 20156 4061 20160
rect 3997 20100 4001 20156
rect 4001 20100 4057 20156
rect 4057 20100 4061 20156
rect 3997 20096 4061 20100
rect 4077 20156 4141 20160
rect 4077 20100 4081 20156
rect 4081 20100 4137 20156
rect 4137 20100 4141 20156
rect 4077 20096 4141 20100
rect 4157 20156 4221 20160
rect 4157 20100 4161 20156
rect 4161 20100 4217 20156
rect 4217 20100 4221 20156
rect 4157 20096 4221 20100
rect 9848 20156 9912 20160
rect 9848 20100 9852 20156
rect 9852 20100 9908 20156
rect 9908 20100 9912 20156
rect 9848 20096 9912 20100
rect 9928 20156 9992 20160
rect 9928 20100 9932 20156
rect 9932 20100 9988 20156
rect 9988 20100 9992 20156
rect 9928 20096 9992 20100
rect 10008 20156 10072 20160
rect 10008 20100 10012 20156
rect 10012 20100 10068 20156
rect 10068 20100 10072 20156
rect 10008 20096 10072 20100
rect 10088 20156 10152 20160
rect 10088 20100 10092 20156
rect 10092 20100 10148 20156
rect 10148 20100 10152 20156
rect 10088 20096 10152 20100
rect 15778 20156 15842 20160
rect 15778 20100 15782 20156
rect 15782 20100 15838 20156
rect 15838 20100 15842 20156
rect 15778 20096 15842 20100
rect 15858 20156 15922 20160
rect 15858 20100 15862 20156
rect 15862 20100 15918 20156
rect 15918 20100 15922 20156
rect 15858 20096 15922 20100
rect 15938 20156 16002 20160
rect 15938 20100 15942 20156
rect 15942 20100 15998 20156
rect 15998 20100 16002 20156
rect 15938 20096 16002 20100
rect 16018 20156 16082 20160
rect 16018 20100 16022 20156
rect 16022 20100 16078 20156
rect 16078 20100 16082 20156
rect 16018 20096 16082 20100
rect 6882 19612 6946 19616
rect 6882 19556 6886 19612
rect 6886 19556 6942 19612
rect 6942 19556 6946 19612
rect 6882 19552 6946 19556
rect 6962 19612 7026 19616
rect 6962 19556 6966 19612
rect 6966 19556 7022 19612
rect 7022 19556 7026 19612
rect 6962 19552 7026 19556
rect 7042 19612 7106 19616
rect 7042 19556 7046 19612
rect 7046 19556 7102 19612
rect 7102 19556 7106 19612
rect 7042 19552 7106 19556
rect 7122 19612 7186 19616
rect 7122 19556 7126 19612
rect 7126 19556 7182 19612
rect 7182 19556 7186 19612
rect 7122 19552 7186 19556
rect 12813 19612 12877 19616
rect 12813 19556 12817 19612
rect 12817 19556 12873 19612
rect 12873 19556 12877 19612
rect 12813 19552 12877 19556
rect 12893 19612 12957 19616
rect 12893 19556 12897 19612
rect 12897 19556 12953 19612
rect 12953 19556 12957 19612
rect 12893 19552 12957 19556
rect 12973 19612 13037 19616
rect 12973 19556 12977 19612
rect 12977 19556 13033 19612
rect 13033 19556 13037 19612
rect 12973 19552 13037 19556
rect 13053 19612 13117 19616
rect 13053 19556 13057 19612
rect 13057 19556 13113 19612
rect 13113 19556 13117 19612
rect 13053 19552 13117 19556
rect 3917 19068 3981 19072
rect 3917 19012 3921 19068
rect 3921 19012 3977 19068
rect 3977 19012 3981 19068
rect 3917 19008 3981 19012
rect 3997 19068 4061 19072
rect 3997 19012 4001 19068
rect 4001 19012 4057 19068
rect 4057 19012 4061 19068
rect 3997 19008 4061 19012
rect 4077 19068 4141 19072
rect 4077 19012 4081 19068
rect 4081 19012 4137 19068
rect 4137 19012 4141 19068
rect 4077 19008 4141 19012
rect 4157 19068 4221 19072
rect 4157 19012 4161 19068
rect 4161 19012 4217 19068
rect 4217 19012 4221 19068
rect 4157 19008 4221 19012
rect 9848 19068 9912 19072
rect 9848 19012 9852 19068
rect 9852 19012 9908 19068
rect 9908 19012 9912 19068
rect 9848 19008 9912 19012
rect 9928 19068 9992 19072
rect 9928 19012 9932 19068
rect 9932 19012 9988 19068
rect 9988 19012 9992 19068
rect 9928 19008 9992 19012
rect 10008 19068 10072 19072
rect 10008 19012 10012 19068
rect 10012 19012 10068 19068
rect 10068 19012 10072 19068
rect 10008 19008 10072 19012
rect 10088 19068 10152 19072
rect 10088 19012 10092 19068
rect 10092 19012 10148 19068
rect 10148 19012 10152 19068
rect 10088 19008 10152 19012
rect 15778 19068 15842 19072
rect 15778 19012 15782 19068
rect 15782 19012 15838 19068
rect 15838 19012 15842 19068
rect 15778 19008 15842 19012
rect 15858 19068 15922 19072
rect 15858 19012 15862 19068
rect 15862 19012 15918 19068
rect 15918 19012 15922 19068
rect 15858 19008 15922 19012
rect 15938 19068 16002 19072
rect 15938 19012 15942 19068
rect 15942 19012 15998 19068
rect 15998 19012 16002 19068
rect 15938 19008 16002 19012
rect 16018 19068 16082 19072
rect 16018 19012 16022 19068
rect 16022 19012 16078 19068
rect 16078 19012 16082 19068
rect 16018 19008 16082 19012
rect 6882 18524 6946 18528
rect 6882 18468 6886 18524
rect 6886 18468 6942 18524
rect 6942 18468 6946 18524
rect 6882 18464 6946 18468
rect 6962 18524 7026 18528
rect 6962 18468 6966 18524
rect 6966 18468 7022 18524
rect 7022 18468 7026 18524
rect 6962 18464 7026 18468
rect 7042 18524 7106 18528
rect 7042 18468 7046 18524
rect 7046 18468 7102 18524
rect 7102 18468 7106 18524
rect 7042 18464 7106 18468
rect 7122 18524 7186 18528
rect 7122 18468 7126 18524
rect 7126 18468 7182 18524
rect 7182 18468 7186 18524
rect 7122 18464 7186 18468
rect 12813 18524 12877 18528
rect 12813 18468 12817 18524
rect 12817 18468 12873 18524
rect 12873 18468 12877 18524
rect 12813 18464 12877 18468
rect 12893 18524 12957 18528
rect 12893 18468 12897 18524
rect 12897 18468 12953 18524
rect 12953 18468 12957 18524
rect 12893 18464 12957 18468
rect 12973 18524 13037 18528
rect 12973 18468 12977 18524
rect 12977 18468 13033 18524
rect 13033 18468 13037 18524
rect 12973 18464 13037 18468
rect 13053 18524 13117 18528
rect 13053 18468 13057 18524
rect 13057 18468 13113 18524
rect 13113 18468 13117 18524
rect 13053 18464 13117 18468
rect 3917 17980 3981 17984
rect 3917 17924 3921 17980
rect 3921 17924 3977 17980
rect 3977 17924 3981 17980
rect 3917 17920 3981 17924
rect 3997 17980 4061 17984
rect 3997 17924 4001 17980
rect 4001 17924 4057 17980
rect 4057 17924 4061 17980
rect 3997 17920 4061 17924
rect 4077 17980 4141 17984
rect 4077 17924 4081 17980
rect 4081 17924 4137 17980
rect 4137 17924 4141 17980
rect 4077 17920 4141 17924
rect 4157 17980 4221 17984
rect 4157 17924 4161 17980
rect 4161 17924 4217 17980
rect 4217 17924 4221 17980
rect 4157 17920 4221 17924
rect 9848 17980 9912 17984
rect 9848 17924 9852 17980
rect 9852 17924 9908 17980
rect 9908 17924 9912 17980
rect 9848 17920 9912 17924
rect 9928 17980 9992 17984
rect 9928 17924 9932 17980
rect 9932 17924 9988 17980
rect 9988 17924 9992 17980
rect 9928 17920 9992 17924
rect 10008 17980 10072 17984
rect 10008 17924 10012 17980
rect 10012 17924 10068 17980
rect 10068 17924 10072 17980
rect 10008 17920 10072 17924
rect 10088 17980 10152 17984
rect 10088 17924 10092 17980
rect 10092 17924 10148 17980
rect 10148 17924 10152 17980
rect 10088 17920 10152 17924
rect 15778 17980 15842 17984
rect 15778 17924 15782 17980
rect 15782 17924 15838 17980
rect 15838 17924 15842 17980
rect 15778 17920 15842 17924
rect 15858 17980 15922 17984
rect 15858 17924 15862 17980
rect 15862 17924 15918 17980
rect 15918 17924 15922 17980
rect 15858 17920 15922 17924
rect 15938 17980 16002 17984
rect 15938 17924 15942 17980
rect 15942 17924 15998 17980
rect 15998 17924 16002 17980
rect 15938 17920 16002 17924
rect 16018 17980 16082 17984
rect 16018 17924 16022 17980
rect 16022 17924 16078 17980
rect 16078 17924 16082 17980
rect 16018 17920 16082 17924
rect 6882 17436 6946 17440
rect 6882 17380 6886 17436
rect 6886 17380 6942 17436
rect 6942 17380 6946 17436
rect 6882 17376 6946 17380
rect 6962 17436 7026 17440
rect 6962 17380 6966 17436
rect 6966 17380 7022 17436
rect 7022 17380 7026 17436
rect 6962 17376 7026 17380
rect 7042 17436 7106 17440
rect 7042 17380 7046 17436
rect 7046 17380 7102 17436
rect 7102 17380 7106 17436
rect 7042 17376 7106 17380
rect 7122 17436 7186 17440
rect 7122 17380 7126 17436
rect 7126 17380 7182 17436
rect 7182 17380 7186 17436
rect 7122 17376 7186 17380
rect 12813 17436 12877 17440
rect 12813 17380 12817 17436
rect 12817 17380 12873 17436
rect 12873 17380 12877 17436
rect 12813 17376 12877 17380
rect 12893 17436 12957 17440
rect 12893 17380 12897 17436
rect 12897 17380 12953 17436
rect 12953 17380 12957 17436
rect 12893 17376 12957 17380
rect 12973 17436 13037 17440
rect 12973 17380 12977 17436
rect 12977 17380 13033 17436
rect 13033 17380 13037 17436
rect 12973 17376 13037 17380
rect 13053 17436 13117 17440
rect 13053 17380 13057 17436
rect 13057 17380 13113 17436
rect 13113 17380 13117 17436
rect 13053 17376 13117 17380
rect 3917 16892 3981 16896
rect 3917 16836 3921 16892
rect 3921 16836 3977 16892
rect 3977 16836 3981 16892
rect 3917 16832 3981 16836
rect 3997 16892 4061 16896
rect 3997 16836 4001 16892
rect 4001 16836 4057 16892
rect 4057 16836 4061 16892
rect 3997 16832 4061 16836
rect 4077 16892 4141 16896
rect 4077 16836 4081 16892
rect 4081 16836 4137 16892
rect 4137 16836 4141 16892
rect 4077 16832 4141 16836
rect 4157 16892 4221 16896
rect 4157 16836 4161 16892
rect 4161 16836 4217 16892
rect 4217 16836 4221 16892
rect 4157 16832 4221 16836
rect 9848 16892 9912 16896
rect 9848 16836 9852 16892
rect 9852 16836 9908 16892
rect 9908 16836 9912 16892
rect 9848 16832 9912 16836
rect 9928 16892 9992 16896
rect 9928 16836 9932 16892
rect 9932 16836 9988 16892
rect 9988 16836 9992 16892
rect 9928 16832 9992 16836
rect 10008 16892 10072 16896
rect 10008 16836 10012 16892
rect 10012 16836 10068 16892
rect 10068 16836 10072 16892
rect 10008 16832 10072 16836
rect 10088 16892 10152 16896
rect 10088 16836 10092 16892
rect 10092 16836 10148 16892
rect 10148 16836 10152 16892
rect 10088 16832 10152 16836
rect 15778 16892 15842 16896
rect 15778 16836 15782 16892
rect 15782 16836 15838 16892
rect 15838 16836 15842 16892
rect 15778 16832 15842 16836
rect 15858 16892 15922 16896
rect 15858 16836 15862 16892
rect 15862 16836 15918 16892
rect 15918 16836 15922 16892
rect 15858 16832 15922 16836
rect 15938 16892 16002 16896
rect 15938 16836 15942 16892
rect 15942 16836 15998 16892
rect 15998 16836 16002 16892
rect 15938 16832 16002 16836
rect 16018 16892 16082 16896
rect 16018 16836 16022 16892
rect 16022 16836 16078 16892
rect 16078 16836 16082 16892
rect 16018 16832 16082 16836
rect 6882 16348 6946 16352
rect 6882 16292 6886 16348
rect 6886 16292 6942 16348
rect 6942 16292 6946 16348
rect 6882 16288 6946 16292
rect 6962 16348 7026 16352
rect 6962 16292 6966 16348
rect 6966 16292 7022 16348
rect 7022 16292 7026 16348
rect 6962 16288 7026 16292
rect 7042 16348 7106 16352
rect 7042 16292 7046 16348
rect 7046 16292 7102 16348
rect 7102 16292 7106 16348
rect 7042 16288 7106 16292
rect 7122 16348 7186 16352
rect 7122 16292 7126 16348
rect 7126 16292 7182 16348
rect 7182 16292 7186 16348
rect 7122 16288 7186 16292
rect 12813 16348 12877 16352
rect 12813 16292 12817 16348
rect 12817 16292 12873 16348
rect 12873 16292 12877 16348
rect 12813 16288 12877 16292
rect 12893 16348 12957 16352
rect 12893 16292 12897 16348
rect 12897 16292 12953 16348
rect 12953 16292 12957 16348
rect 12893 16288 12957 16292
rect 12973 16348 13037 16352
rect 12973 16292 12977 16348
rect 12977 16292 13033 16348
rect 13033 16292 13037 16348
rect 12973 16288 13037 16292
rect 13053 16348 13117 16352
rect 13053 16292 13057 16348
rect 13057 16292 13113 16348
rect 13113 16292 13117 16348
rect 13053 16288 13117 16292
rect 3917 15804 3981 15808
rect 3917 15748 3921 15804
rect 3921 15748 3977 15804
rect 3977 15748 3981 15804
rect 3917 15744 3981 15748
rect 3997 15804 4061 15808
rect 3997 15748 4001 15804
rect 4001 15748 4057 15804
rect 4057 15748 4061 15804
rect 3997 15744 4061 15748
rect 4077 15804 4141 15808
rect 4077 15748 4081 15804
rect 4081 15748 4137 15804
rect 4137 15748 4141 15804
rect 4077 15744 4141 15748
rect 4157 15804 4221 15808
rect 4157 15748 4161 15804
rect 4161 15748 4217 15804
rect 4217 15748 4221 15804
rect 4157 15744 4221 15748
rect 9848 15804 9912 15808
rect 9848 15748 9852 15804
rect 9852 15748 9908 15804
rect 9908 15748 9912 15804
rect 9848 15744 9912 15748
rect 9928 15804 9992 15808
rect 9928 15748 9932 15804
rect 9932 15748 9988 15804
rect 9988 15748 9992 15804
rect 9928 15744 9992 15748
rect 10008 15804 10072 15808
rect 10008 15748 10012 15804
rect 10012 15748 10068 15804
rect 10068 15748 10072 15804
rect 10008 15744 10072 15748
rect 10088 15804 10152 15808
rect 10088 15748 10092 15804
rect 10092 15748 10148 15804
rect 10148 15748 10152 15804
rect 10088 15744 10152 15748
rect 15778 15804 15842 15808
rect 15778 15748 15782 15804
rect 15782 15748 15838 15804
rect 15838 15748 15842 15804
rect 15778 15744 15842 15748
rect 15858 15804 15922 15808
rect 15858 15748 15862 15804
rect 15862 15748 15918 15804
rect 15918 15748 15922 15804
rect 15858 15744 15922 15748
rect 15938 15804 16002 15808
rect 15938 15748 15942 15804
rect 15942 15748 15998 15804
rect 15998 15748 16002 15804
rect 15938 15744 16002 15748
rect 16018 15804 16082 15808
rect 16018 15748 16022 15804
rect 16022 15748 16078 15804
rect 16078 15748 16082 15804
rect 16018 15744 16082 15748
rect 6882 15260 6946 15264
rect 6882 15204 6886 15260
rect 6886 15204 6942 15260
rect 6942 15204 6946 15260
rect 6882 15200 6946 15204
rect 6962 15260 7026 15264
rect 6962 15204 6966 15260
rect 6966 15204 7022 15260
rect 7022 15204 7026 15260
rect 6962 15200 7026 15204
rect 7042 15260 7106 15264
rect 7042 15204 7046 15260
rect 7046 15204 7102 15260
rect 7102 15204 7106 15260
rect 7042 15200 7106 15204
rect 7122 15260 7186 15264
rect 7122 15204 7126 15260
rect 7126 15204 7182 15260
rect 7182 15204 7186 15260
rect 7122 15200 7186 15204
rect 12813 15260 12877 15264
rect 12813 15204 12817 15260
rect 12817 15204 12873 15260
rect 12873 15204 12877 15260
rect 12813 15200 12877 15204
rect 12893 15260 12957 15264
rect 12893 15204 12897 15260
rect 12897 15204 12953 15260
rect 12953 15204 12957 15260
rect 12893 15200 12957 15204
rect 12973 15260 13037 15264
rect 12973 15204 12977 15260
rect 12977 15204 13033 15260
rect 13033 15204 13037 15260
rect 12973 15200 13037 15204
rect 13053 15260 13117 15264
rect 13053 15204 13057 15260
rect 13057 15204 13113 15260
rect 13113 15204 13117 15260
rect 13053 15200 13117 15204
rect 3917 14716 3981 14720
rect 3917 14660 3921 14716
rect 3921 14660 3977 14716
rect 3977 14660 3981 14716
rect 3917 14656 3981 14660
rect 3997 14716 4061 14720
rect 3997 14660 4001 14716
rect 4001 14660 4057 14716
rect 4057 14660 4061 14716
rect 3997 14656 4061 14660
rect 4077 14716 4141 14720
rect 4077 14660 4081 14716
rect 4081 14660 4137 14716
rect 4137 14660 4141 14716
rect 4077 14656 4141 14660
rect 4157 14716 4221 14720
rect 4157 14660 4161 14716
rect 4161 14660 4217 14716
rect 4217 14660 4221 14716
rect 4157 14656 4221 14660
rect 9848 14716 9912 14720
rect 9848 14660 9852 14716
rect 9852 14660 9908 14716
rect 9908 14660 9912 14716
rect 9848 14656 9912 14660
rect 9928 14716 9992 14720
rect 9928 14660 9932 14716
rect 9932 14660 9988 14716
rect 9988 14660 9992 14716
rect 9928 14656 9992 14660
rect 10008 14716 10072 14720
rect 10008 14660 10012 14716
rect 10012 14660 10068 14716
rect 10068 14660 10072 14716
rect 10008 14656 10072 14660
rect 10088 14716 10152 14720
rect 10088 14660 10092 14716
rect 10092 14660 10148 14716
rect 10148 14660 10152 14716
rect 10088 14656 10152 14660
rect 15778 14716 15842 14720
rect 15778 14660 15782 14716
rect 15782 14660 15838 14716
rect 15838 14660 15842 14716
rect 15778 14656 15842 14660
rect 15858 14716 15922 14720
rect 15858 14660 15862 14716
rect 15862 14660 15918 14716
rect 15918 14660 15922 14716
rect 15858 14656 15922 14660
rect 15938 14716 16002 14720
rect 15938 14660 15942 14716
rect 15942 14660 15998 14716
rect 15998 14660 16002 14716
rect 15938 14656 16002 14660
rect 16018 14716 16082 14720
rect 16018 14660 16022 14716
rect 16022 14660 16078 14716
rect 16078 14660 16082 14716
rect 16018 14656 16082 14660
rect 6882 14172 6946 14176
rect 6882 14116 6886 14172
rect 6886 14116 6942 14172
rect 6942 14116 6946 14172
rect 6882 14112 6946 14116
rect 6962 14172 7026 14176
rect 6962 14116 6966 14172
rect 6966 14116 7022 14172
rect 7022 14116 7026 14172
rect 6962 14112 7026 14116
rect 7042 14172 7106 14176
rect 7042 14116 7046 14172
rect 7046 14116 7102 14172
rect 7102 14116 7106 14172
rect 7042 14112 7106 14116
rect 7122 14172 7186 14176
rect 7122 14116 7126 14172
rect 7126 14116 7182 14172
rect 7182 14116 7186 14172
rect 7122 14112 7186 14116
rect 12813 14172 12877 14176
rect 12813 14116 12817 14172
rect 12817 14116 12873 14172
rect 12873 14116 12877 14172
rect 12813 14112 12877 14116
rect 12893 14172 12957 14176
rect 12893 14116 12897 14172
rect 12897 14116 12953 14172
rect 12953 14116 12957 14172
rect 12893 14112 12957 14116
rect 12973 14172 13037 14176
rect 12973 14116 12977 14172
rect 12977 14116 13033 14172
rect 13033 14116 13037 14172
rect 12973 14112 13037 14116
rect 13053 14172 13117 14176
rect 13053 14116 13057 14172
rect 13057 14116 13113 14172
rect 13113 14116 13117 14172
rect 13053 14112 13117 14116
rect 3917 13628 3981 13632
rect 3917 13572 3921 13628
rect 3921 13572 3977 13628
rect 3977 13572 3981 13628
rect 3917 13568 3981 13572
rect 3997 13628 4061 13632
rect 3997 13572 4001 13628
rect 4001 13572 4057 13628
rect 4057 13572 4061 13628
rect 3997 13568 4061 13572
rect 4077 13628 4141 13632
rect 4077 13572 4081 13628
rect 4081 13572 4137 13628
rect 4137 13572 4141 13628
rect 4077 13568 4141 13572
rect 4157 13628 4221 13632
rect 4157 13572 4161 13628
rect 4161 13572 4217 13628
rect 4217 13572 4221 13628
rect 4157 13568 4221 13572
rect 9848 13628 9912 13632
rect 9848 13572 9852 13628
rect 9852 13572 9908 13628
rect 9908 13572 9912 13628
rect 9848 13568 9912 13572
rect 9928 13628 9992 13632
rect 9928 13572 9932 13628
rect 9932 13572 9988 13628
rect 9988 13572 9992 13628
rect 9928 13568 9992 13572
rect 10008 13628 10072 13632
rect 10008 13572 10012 13628
rect 10012 13572 10068 13628
rect 10068 13572 10072 13628
rect 10008 13568 10072 13572
rect 10088 13628 10152 13632
rect 10088 13572 10092 13628
rect 10092 13572 10148 13628
rect 10148 13572 10152 13628
rect 10088 13568 10152 13572
rect 15778 13628 15842 13632
rect 15778 13572 15782 13628
rect 15782 13572 15838 13628
rect 15838 13572 15842 13628
rect 15778 13568 15842 13572
rect 15858 13628 15922 13632
rect 15858 13572 15862 13628
rect 15862 13572 15918 13628
rect 15918 13572 15922 13628
rect 15858 13568 15922 13572
rect 15938 13628 16002 13632
rect 15938 13572 15942 13628
rect 15942 13572 15998 13628
rect 15998 13572 16002 13628
rect 15938 13568 16002 13572
rect 16018 13628 16082 13632
rect 16018 13572 16022 13628
rect 16022 13572 16078 13628
rect 16078 13572 16082 13628
rect 16018 13568 16082 13572
rect 6882 13084 6946 13088
rect 6882 13028 6886 13084
rect 6886 13028 6942 13084
rect 6942 13028 6946 13084
rect 6882 13024 6946 13028
rect 6962 13084 7026 13088
rect 6962 13028 6966 13084
rect 6966 13028 7022 13084
rect 7022 13028 7026 13084
rect 6962 13024 7026 13028
rect 7042 13084 7106 13088
rect 7042 13028 7046 13084
rect 7046 13028 7102 13084
rect 7102 13028 7106 13084
rect 7042 13024 7106 13028
rect 7122 13084 7186 13088
rect 7122 13028 7126 13084
rect 7126 13028 7182 13084
rect 7182 13028 7186 13084
rect 7122 13024 7186 13028
rect 12813 13084 12877 13088
rect 12813 13028 12817 13084
rect 12817 13028 12873 13084
rect 12873 13028 12877 13084
rect 12813 13024 12877 13028
rect 12893 13084 12957 13088
rect 12893 13028 12897 13084
rect 12897 13028 12953 13084
rect 12953 13028 12957 13084
rect 12893 13024 12957 13028
rect 12973 13084 13037 13088
rect 12973 13028 12977 13084
rect 12977 13028 13033 13084
rect 13033 13028 13037 13084
rect 12973 13024 13037 13028
rect 13053 13084 13117 13088
rect 13053 13028 13057 13084
rect 13057 13028 13113 13084
rect 13113 13028 13117 13084
rect 13053 13024 13117 13028
rect 3917 12540 3981 12544
rect 3917 12484 3921 12540
rect 3921 12484 3977 12540
rect 3977 12484 3981 12540
rect 3917 12480 3981 12484
rect 3997 12540 4061 12544
rect 3997 12484 4001 12540
rect 4001 12484 4057 12540
rect 4057 12484 4061 12540
rect 3997 12480 4061 12484
rect 4077 12540 4141 12544
rect 4077 12484 4081 12540
rect 4081 12484 4137 12540
rect 4137 12484 4141 12540
rect 4077 12480 4141 12484
rect 4157 12540 4221 12544
rect 4157 12484 4161 12540
rect 4161 12484 4217 12540
rect 4217 12484 4221 12540
rect 4157 12480 4221 12484
rect 9848 12540 9912 12544
rect 9848 12484 9852 12540
rect 9852 12484 9908 12540
rect 9908 12484 9912 12540
rect 9848 12480 9912 12484
rect 9928 12540 9992 12544
rect 9928 12484 9932 12540
rect 9932 12484 9988 12540
rect 9988 12484 9992 12540
rect 9928 12480 9992 12484
rect 10008 12540 10072 12544
rect 10008 12484 10012 12540
rect 10012 12484 10068 12540
rect 10068 12484 10072 12540
rect 10008 12480 10072 12484
rect 10088 12540 10152 12544
rect 10088 12484 10092 12540
rect 10092 12484 10148 12540
rect 10148 12484 10152 12540
rect 10088 12480 10152 12484
rect 15778 12540 15842 12544
rect 15778 12484 15782 12540
rect 15782 12484 15838 12540
rect 15838 12484 15842 12540
rect 15778 12480 15842 12484
rect 15858 12540 15922 12544
rect 15858 12484 15862 12540
rect 15862 12484 15918 12540
rect 15918 12484 15922 12540
rect 15858 12480 15922 12484
rect 15938 12540 16002 12544
rect 15938 12484 15942 12540
rect 15942 12484 15998 12540
rect 15998 12484 16002 12540
rect 15938 12480 16002 12484
rect 16018 12540 16082 12544
rect 16018 12484 16022 12540
rect 16022 12484 16078 12540
rect 16078 12484 16082 12540
rect 16018 12480 16082 12484
rect 6882 11996 6946 12000
rect 6882 11940 6886 11996
rect 6886 11940 6942 11996
rect 6942 11940 6946 11996
rect 6882 11936 6946 11940
rect 6962 11996 7026 12000
rect 6962 11940 6966 11996
rect 6966 11940 7022 11996
rect 7022 11940 7026 11996
rect 6962 11936 7026 11940
rect 7042 11996 7106 12000
rect 7042 11940 7046 11996
rect 7046 11940 7102 11996
rect 7102 11940 7106 11996
rect 7042 11936 7106 11940
rect 7122 11996 7186 12000
rect 7122 11940 7126 11996
rect 7126 11940 7182 11996
rect 7182 11940 7186 11996
rect 7122 11936 7186 11940
rect 12813 11996 12877 12000
rect 12813 11940 12817 11996
rect 12817 11940 12873 11996
rect 12873 11940 12877 11996
rect 12813 11936 12877 11940
rect 12893 11996 12957 12000
rect 12893 11940 12897 11996
rect 12897 11940 12953 11996
rect 12953 11940 12957 11996
rect 12893 11936 12957 11940
rect 12973 11996 13037 12000
rect 12973 11940 12977 11996
rect 12977 11940 13033 11996
rect 13033 11940 13037 11996
rect 12973 11936 13037 11940
rect 13053 11996 13117 12000
rect 13053 11940 13057 11996
rect 13057 11940 13113 11996
rect 13113 11940 13117 11996
rect 13053 11936 13117 11940
rect 3917 11452 3981 11456
rect 3917 11396 3921 11452
rect 3921 11396 3977 11452
rect 3977 11396 3981 11452
rect 3917 11392 3981 11396
rect 3997 11452 4061 11456
rect 3997 11396 4001 11452
rect 4001 11396 4057 11452
rect 4057 11396 4061 11452
rect 3997 11392 4061 11396
rect 4077 11452 4141 11456
rect 4077 11396 4081 11452
rect 4081 11396 4137 11452
rect 4137 11396 4141 11452
rect 4077 11392 4141 11396
rect 4157 11452 4221 11456
rect 4157 11396 4161 11452
rect 4161 11396 4217 11452
rect 4217 11396 4221 11452
rect 4157 11392 4221 11396
rect 9848 11452 9912 11456
rect 9848 11396 9852 11452
rect 9852 11396 9908 11452
rect 9908 11396 9912 11452
rect 9848 11392 9912 11396
rect 9928 11452 9992 11456
rect 9928 11396 9932 11452
rect 9932 11396 9988 11452
rect 9988 11396 9992 11452
rect 9928 11392 9992 11396
rect 10008 11452 10072 11456
rect 10008 11396 10012 11452
rect 10012 11396 10068 11452
rect 10068 11396 10072 11452
rect 10008 11392 10072 11396
rect 10088 11452 10152 11456
rect 10088 11396 10092 11452
rect 10092 11396 10148 11452
rect 10148 11396 10152 11452
rect 10088 11392 10152 11396
rect 15778 11452 15842 11456
rect 15778 11396 15782 11452
rect 15782 11396 15838 11452
rect 15838 11396 15842 11452
rect 15778 11392 15842 11396
rect 15858 11452 15922 11456
rect 15858 11396 15862 11452
rect 15862 11396 15918 11452
rect 15918 11396 15922 11452
rect 15858 11392 15922 11396
rect 15938 11452 16002 11456
rect 15938 11396 15942 11452
rect 15942 11396 15998 11452
rect 15998 11396 16002 11452
rect 15938 11392 16002 11396
rect 16018 11452 16082 11456
rect 16018 11396 16022 11452
rect 16022 11396 16078 11452
rect 16078 11396 16082 11452
rect 16018 11392 16082 11396
rect 6882 10908 6946 10912
rect 6882 10852 6886 10908
rect 6886 10852 6942 10908
rect 6942 10852 6946 10908
rect 6882 10848 6946 10852
rect 6962 10908 7026 10912
rect 6962 10852 6966 10908
rect 6966 10852 7022 10908
rect 7022 10852 7026 10908
rect 6962 10848 7026 10852
rect 7042 10908 7106 10912
rect 7042 10852 7046 10908
rect 7046 10852 7102 10908
rect 7102 10852 7106 10908
rect 7042 10848 7106 10852
rect 7122 10908 7186 10912
rect 7122 10852 7126 10908
rect 7126 10852 7182 10908
rect 7182 10852 7186 10908
rect 7122 10848 7186 10852
rect 12813 10908 12877 10912
rect 12813 10852 12817 10908
rect 12817 10852 12873 10908
rect 12873 10852 12877 10908
rect 12813 10848 12877 10852
rect 12893 10908 12957 10912
rect 12893 10852 12897 10908
rect 12897 10852 12953 10908
rect 12953 10852 12957 10908
rect 12893 10848 12957 10852
rect 12973 10908 13037 10912
rect 12973 10852 12977 10908
rect 12977 10852 13033 10908
rect 13033 10852 13037 10908
rect 12973 10848 13037 10852
rect 13053 10908 13117 10912
rect 13053 10852 13057 10908
rect 13057 10852 13113 10908
rect 13113 10852 13117 10908
rect 13053 10848 13117 10852
rect 3917 10364 3981 10368
rect 3917 10308 3921 10364
rect 3921 10308 3977 10364
rect 3977 10308 3981 10364
rect 3917 10304 3981 10308
rect 3997 10364 4061 10368
rect 3997 10308 4001 10364
rect 4001 10308 4057 10364
rect 4057 10308 4061 10364
rect 3997 10304 4061 10308
rect 4077 10364 4141 10368
rect 4077 10308 4081 10364
rect 4081 10308 4137 10364
rect 4137 10308 4141 10364
rect 4077 10304 4141 10308
rect 4157 10364 4221 10368
rect 4157 10308 4161 10364
rect 4161 10308 4217 10364
rect 4217 10308 4221 10364
rect 4157 10304 4221 10308
rect 9848 10364 9912 10368
rect 9848 10308 9852 10364
rect 9852 10308 9908 10364
rect 9908 10308 9912 10364
rect 9848 10304 9912 10308
rect 9928 10364 9992 10368
rect 9928 10308 9932 10364
rect 9932 10308 9988 10364
rect 9988 10308 9992 10364
rect 9928 10304 9992 10308
rect 10008 10364 10072 10368
rect 10008 10308 10012 10364
rect 10012 10308 10068 10364
rect 10068 10308 10072 10364
rect 10008 10304 10072 10308
rect 10088 10364 10152 10368
rect 10088 10308 10092 10364
rect 10092 10308 10148 10364
rect 10148 10308 10152 10364
rect 10088 10304 10152 10308
rect 15778 10364 15842 10368
rect 15778 10308 15782 10364
rect 15782 10308 15838 10364
rect 15838 10308 15842 10364
rect 15778 10304 15842 10308
rect 15858 10364 15922 10368
rect 15858 10308 15862 10364
rect 15862 10308 15918 10364
rect 15918 10308 15922 10364
rect 15858 10304 15922 10308
rect 15938 10364 16002 10368
rect 15938 10308 15942 10364
rect 15942 10308 15998 10364
rect 15998 10308 16002 10364
rect 15938 10304 16002 10308
rect 16018 10364 16082 10368
rect 16018 10308 16022 10364
rect 16022 10308 16078 10364
rect 16078 10308 16082 10364
rect 16018 10304 16082 10308
rect 6882 9820 6946 9824
rect 6882 9764 6886 9820
rect 6886 9764 6942 9820
rect 6942 9764 6946 9820
rect 6882 9760 6946 9764
rect 6962 9820 7026 9824
rect 6962 9764 6966 9820
rect 6966 9764 7022 9820
rect 7022 9764 7026 9820
rect 6962 9760 7026 9764
rect 7042 9820 7106 9824
rect 7042 9764 7046 9820
rect 7046 9764 7102 9820
rect 7102 9764 7106 9820
rect 7042 9760 7106 9764
rect 7122 9820 7186 9824
rect 7122 9764 7126 9820
rect 7126 9764 7182 9820
rect 7182 9764 7186 9820
rect 7122 9760 7186 9764
rect 12813 9820 12877 9824
rect 12813 9764 12817 9820
rect 12817 9764 12873 9820
rect 12873 9764 12877 9820
rect 12813 9760 12877 9764
rect 12893 9820 12957 9824
rect 12893 9764 12897 9820
rect 12897 9764 12953 9820
rect 12953 9764 12957 9820
rect 12893 9760 12957 9764
rect 12973 9820 13037 9824
rect 12973 9764 12977 9820
rect 12977 9764 13033 9820
rect 13033 9764 13037 9820
rect 12973 9760 13037 9764
rect 13053 9820 13117 9824
rect 13053 9764 13057 9820
rect 13057 9764 13113 9820
rect 13113 9764 13117 9820
rect 13053 9760 13117 9764
rect 3917 9276 3981 9280
rect 3917 9220 3921 9276
rect 3921 9220 3977 9276
rect 3977 9220 3981 9276
rect 3917 9216 3981 9220
rect 3997 9276 4061 9280
rect 3997 9220 4001 9276
rect 4001 9220 4057 9276
rect 4057 9220 4061 9276
rect 3997 9216 4061 9220
rect 4077 9276 4141 9280
rect 4077 9220 4081 9276
rect 4081 9220 4137 9276
rect 4137 9220 4141 9276
rect 4077 9216 4141 9220
rect 4157 9276 4221 9280
rect 4157 9220 4161 9276
rect 4161 9220 4217 9276
rect 4217 9220 4221 9276
rect 4157 9216 4221 9220
rect 9848 9276 9912 9280
rect 9848 9220 9852 9276
rect 9852 9220 9908 9276
rect 9908 9220 9912 9276
rect 9848 9216 9912 9220
rect 9928 9276 9992 9280
rect 9928 9220 9932 9276
rect 9932 9220 9988 9276
rect 9988 9220 9992 9276
rect 9928 9216 9992 9220
rect 10008 9276 10072 9280
rect 10008 9220 10012 9276
rect 10012 9220 10068 9276
rect 10068 9220 10072 9276
rect 10008 9216 10072 9220
rect 10088 9276 10152 9280
rect 10088 9220 10092 9276
rect 10092 9220 10148 9276
rect 10148 9220 10152 9276
rect 10088 9216 10152 9220
rect 15778 9276 15842 9280
rect 15778 9220 15782 9276
rect 15782 9220 15838 9276
rect 15838 9220 15842 9276
rect 15778 9216 15842 9220
rect 15858 9276 15922 9280
rect 15858 9220 15862 9276
rect 15862 9220 15918 9276
rect 15918 9220 15922 9276
rect 15858 9216 15922 9220
rect 15938 9276 16002 9280
rect 15938 9220 15942 9276
rect 15942 9220 15998 9276
rect 15998 9220 16002 9276
rect 15938 9216 16002 9220
rect 16018 9276 16082 9280
rect 16018 9220 16022 9276
rect 16022 9220 16078 9276
rect 16078 9220 16082 9276
rect 16018 9216 16082 9220
rect 6882 8732 6946 8736
rect 6882 8676 6886 8732
rect 6886 8676 6942 8732
rect 6942 8676 6946 8732
rect 6882 8672 6946 8676
rect 6962 8732 7026 8736
rect 6962 8676 6966 8732
rect 6966 8676 7022 8732
rect 7022 8676 7026 8732
rect 6962 8672 7026 8676
rect 7042 8732 7106 8736
rect 7042 8676 7046 8732
rect 7046 8676 7102 8732
rect 7102 8676 7106 8732
rect 7042 8672 7106 8676
rect 7122 8732 7186 8736
rect 7122 8676 7126 8732
rect 7126 8676 7182 8732
rect 7182 8676 7186 8732
rect 7122 8672 7186 8676
rect 12813 8732 12877 8736
rect 12813 8676 12817 8732
rect 12817 8676 12873 8732
rect 12873 8676 12877 8732
rect 12813 8672 12877 8676
rect 12893 8732 12957 8736
rect 12893 8676 12897 8732
rect 12897 8676 12953 8732
rect 12953 8676 12957 8732
rect 12893 8672 12957 8676
rect 12973 8732 13037 8736
rect 12973 8676 12977 8732
rect 12977 8676 13033 8732
rect 13033 8676 13037 8732
rect 12973 8672 13037 8676
rect 13053 8732 13117 8736
rect 13053 8676 13057 8732
rect 13057 8676 13113 8732
rect 13113 8676 13117 8732
rect 13053 8672 13117 8676
rect 3917 8188 3981 8192
rect 3917 8132 3921 8188
rect 3921 8132 3977 8188
rect 3977 8132 3981 8188
rect 3917 8128 3981 8132
rect 3997 8188 4061 8192
rect 3997 8132 4001 8188
rect 4001 8132 4057 8188
rect 4057 8132 4061 8188
rect 3997 8128 4061 8132
rect 4077 8188 4141 8192
rect 4077 8132 4081 8188
rect 4081 8132 4137 8188
rect 4137 8132 4141 8188
rect 4077 8128 4141 8132
rect 4157 8188 4221 8192
rect 4157 8132 4161 8188
rect 4161 8132 4217 8188
rect 4217 8132 4221 8188
rect 4157 8128 4221 8132
rect 9848 8188 9912 8192
rect 9848 8132 9852 8188
rect 9852 8132 9908 8188
rect 9908 8132 9912 8188
rect 9848 8128 9912 8132
rect 9928 8188 9992 8192
rect 9928 8132 9932 8188
rect 9932 8132 9988 8188
rect 9988 8132 9992 8188
rect 9928 8128 9992 8132
rect 10008 8188 10072 8192
rect 10008 8132 10012 8188
rect 10012 8132 10068 8188
rect 10068 8132 10072 8188
rect 10008 8128 10072 8132
rect 10088 8188 10152 8192
rect 10088 8132 10092 8188
rect 10092 8132 10148 8188
rect 10148 8132 10152 8188
rect 10088 8128 10152 8132
rect 15778 8188 15842 8192
rect 15778 8132 15782 8188
rect 15782 8132 15838 8188
rect 15838 8132 15842 8188
rect 15778 8128 15842 8132
rect 15858 8188 15922 8192
rect 15858 8132 15862 8188
rect 15862 8132 15918 8188
rect 15918 8132 15922 8188
rect 15858 8128 15922 8132
rect 15938 8188 16002 8192
rect 15938 8132 15942 8188
rect 15942 8132 15998 8188
rect 15998 8132 16002 8188
rect 15938 8128 16002 8132
rect 16018 8188 16082 8192
rect 16018 8132 16022 8188
rect 16022 8132 16078 8188
rect 16078 8132 16082 8188
rect 16018 8128 16082 8132
rect 6882 7644 6946 7648
rect 6882 7588 6886 7644
rect 6886 7588 6942 7644
rect 6942 7588 6946 7644
rect 6882 7584 6946 7588
rect 6962 7644 7026 7648
rect 6962 7588 6966 7644
rect 6966 7588 7022 7644
rect 7022 7588 7026 7644
rect 6962 7584 7026 7588
rect 7042 7644 7106 7648
rect 7042 7588 7046 7644
rect 7046 7588 7102 7644
rect 7102 7588 7106 7644
rect 7042 7584 7106 7588
rect 7122 7644 7186 7648
rect 7122 7588 7126 7644
rect 7126 7588 7182 7644
rect 7182 7588 7186 7644
rect 7122 7584 7186 7588
rect 12813 7644 12877 7648
rect 12813 7588 12817 7644
rect 12817 7588 12873 7644
rect 12873 7588 12877 7644
rect 12813 7584 12877 7588
rect 12893 7644 12957 7648
rect 12893 7588 12897 7644
rect 12897 7588 12953 7644
rect 12953 7588 12957 7644
rect 12893 7584 12957 7588
rect 12973 7644 13037 7648
rect 12973 7588 12977 7644
rect 12977 7588 13033 7644
rect 13033 7588 13037 7644
rect 12973 7584 13037 7588
rect 13053 7644 13117 7648
rect 13053 7588 13057 7644
rect 13057 7588 13113 7644
rect 13113 7588 13117 7644
rect 13053 7584 13117 7588
rect 3917 7100 3981 7104
rect 3917 7044 3921 7100
rect 3921 7044 3977 7100
rect 3977 7044 3981 7100
rect 3917 7040 3981 7044
rect 3997 7100 4061 7104
rect 3997 7044 4001 7100
rect 4001 7044 4057 7100
rect 4057 7044 4061 7100
rect 3997 7040 4061 7044
rect 4077 7100 4141 7104
rect 4077 7044 4081 7100
rect 4081 7044 4137 7100
rect 4137 7044 4141 7100
rect 4077 7040 4141 7044
rect 4157 7100 4221 7104
rect 4157 7044 4161 7100
rect 4161 7044 4217 7100
rect 4217 7044 4221 7100
rect 4157 7040 4221 7044
rect 9848 7100 9912 7104
rect 9848 7044 9852 7100
rect 9852 7044 9908 7100
rect 9908 7044 9912 7100
rect 9848 7040 9912 7044
rect 9928 7100 9992 7104
rect 9928 7044 9932 7100
rect 9932 7044 9988 7100
rect 9988 7044 9992 7100
rect 9928 7040 9992 7044
rect 10008 7100 10072 7104
rect 10008 7044 10012 7100
rect 10012 7044 10068 7100
rect 10068 7044 10072 7100
rect 10008 7040 10072 7044
rect 10088 7100 10152 7104
rect 10088 7044 10092 7100
rect 10092 7044 10148 7100
rect 10148 7044 10152 7100
rect 10088 7040 10152 7044
rect 15778 7100 15842 7104
rect 15778 7044 15782 7100
rect 15782 7044 15838 7100
rect 15838 7044 15842 7100
rect 15778 7040 15842 7044
rect 15858 7100 15922 7104
rect 15858 7044 15862 7100
rect 15862 7044 15918 7100
rect 15918 7044 15922 7100
rect 15858 7040 15922 7044
rect 15938 7100 16002 7104
rect 15938 7044 15942 7100
rect 15942 7044 15998 7100
rect 15998 7044 16002 7100
rect 15938 7040 16002 7044
rect 16018 7100 16082 7104
rect 16018 7044 16022 7100
rect 16022 7044 16078 7100
rect 16078 7044 16082 7100
rect 16018 7040 16082 7044
rect 6882 6556 6946 6560
rect 6882 6500 6886 6556
rect 6886 6500 6942 6556
rect 6942 6500 6946 6556
rect 6882 6496 6946 6500
rect 6962 6556 7026 6560
rect 6962 6500 6966 6556
rect 6966 6500 7022 6556
rect 7022 6500 7026 6556
rect 6962 6496 7026 6500
rect 7042 6556 7106 6560
rect 7042 6500 7046 6556
rect 7046 6500 7102 6556
rect 7102 6500 7106 6556
rect 7042 6496 7106 6500
rect 7122 6556 7186 6560
rect 7122 6500 7126 6556
rect 7126 6500 7182 6556
rect 7182 6500 7186 6556
rect 7122 6496 7186 6500
rect 12813 6556 12877 6560
rect 12813 6500 12817 6556
rect 12817 6500 12873 6556
rect 12873 6500 12877 6556
rect 12813 6496 12877 6500
rect 12893 6556 12957 6560
rect 12893 6500 12897 6556
rect 12897 6500 12953 6556
rect 12953 6500 12957 6556
rect 12893 6496 12957 6500
rect 12973 6556 13037 6560
rect 12973 6500 12977 6556
rect 12977 6500 13033 6556
rect 13033 6500 13037 6556
rect 12973 6496 13037 6500
rect 13053 6556 13117 6560
rect 13053 6500 13057 6556
rect 13057 6500 13113 6556
rect 13113 6500 13117 6556
rect 13053 6496 13117 6500
rect 3917 6012 3981 6016
rect 3917 5956 3921 6012
rect 3921 5956 3977 6012
rect 3977 5956 3981 6012
rect 3917 5952 3981 5956
rect 3997 6012 4061 6016
rect 3997 5956 4001 6012
rect 4001 5956 4057 6012
rect 4057 5956 4061 6012
rect 3997 5952 4061 5956
rect 4077 6012 4141 6016
rect 4077 5956 4081 6012
rect 4081 5956 4137 6012
rect 4137 5956 4141 6012
rect 4077 5952 4141 5956
rect 4157 6012 4221 6016
rect 4157 5956 4161 6012
rect 4161 5956 4217 6012
rect 4217 5956 4221 6012
rect 4157 5952 4221 5956
rect 9848 6012 9912 6016
rect 9848 5956 9852 6012
rect 9852 5956 9908 6012
rect 9908 5956 9912 6012
rect 9848 5952 9912 5956
rect 9928 6012 9992 6016
rect 9928 5956 9932 6012
rect 9932 5956 9988 6012
rect 9988 5956 9992 6012
rect 9928 5952 9992 5956
rect 10008 6012 10072 6016
rect 10008 5956 10012 6012
rect 10012 5956 10068 6012
rect 10068 5956 10072 6012
rect 10008 5952 10072 5956
rect 10088 6012 10152 6016
rect 10088 5956 10092 6012
rect 10092 5956 10148 6012
rect 10148 5956 10152 6012
rect 10088 5952 10152 5956
rect 15778 6012 15842 6016
rect 15778 5956 15782 6012
rect 15782 5956 15838 6012
rect 15838 5956 15842 6012
rect 15778 5952 15842 5956
rect 15858 6012 15922 6016
rect 15858 5956 15862 6012
rect 15862 5956 15918 6012
rect 15918 5956 15922 6012
rect 15858 5952 15922 5956
rect 15938 6012 16002 6016
rect 15938 5956 15942 6012
rect 15942 5956 15998 6012
rect 15998 5956 16002 6012
rect 15938 5952 16002 5956
rect 16018 6012 16082 6016
rect 16018 5956 16022 6012
rect 16022 5956 16078 6012
rect 16078 5956 16082 6012
rect 16018 5952 16082 5956
rect 6882 5468 6946 5472
rect 6882 5412 6886 5468
rect 6886 5412 6942 5468
rect 6942 5412 6946 5468
rect 6882 5408 6946 5412
rect 6962 5468 7026 5472
rect 6962 5412 6966 5468
rect 6966 5412 7022 5468
rect 7022 5412 7026 5468
rect 6962 5408 7026 5412
rect 7042 5468 7106 5472
rect 7042 5412 7046 5468
rect 7046 5412 7102 5468
rect 7102 5412 7106 5468
rect 7042 5408 7106 5412
rect 7122 5468 7186 5472
rect 7122 5412 7126 5468
rect 7126 5412 7182 5468
rect 7182 5412 7186 5468
rect 7122 5408 7186 5412
rect 12813 5468 12877 5472
rect 12813 5412 12817 5468
rect 12817 5412 12873 5468
rect 12873 5412 12877 5468
rect 12813 5408 12877 5412
rect 12893 5468 12957 5472
rect 12893 5412 12897 5468
rect 12897 5412 12953 5468
rect 12953 5412 12957 5468
rect 12893 5408 12957 5412
rect 12973 5468 13037 5472
rect 12973 5412 12977 5468
rect 12977 5412 13033 5468
rect 13033 5412 13037 5468
rect 12973 5408 13037 5412
rect 13053 5468 13117 5472
rect 13053 5412 13057 5468
rect 13057 5412 13113 5468
rect 13113 5412 13117 5468
rect 13053 5408 13117 5412
rect 3917 4924 3981 4928
rect 3917 4868 3921 4924
rect 3921 4868 3977 4924
rect 3977 4868 3981 4924
rect 3917 4864 3981 4868
rect 3997 4924 4061 4928
rect 3997 4868 4001 4924
rect 4001 4868 4057 4924
rect 4057 4868 4061 4924
rect 3997 4864 4061 4868
rect 4077 4924 4141 4928
rect 4077 4868 4081 4924
rect 4081 4868 4137 4924
rect 4137 4868 4141 4924
rect 4077 4864 4141 4868
rect 4157 4924 4221 4928
rect 4157 4868 4161 4924
rect 4161 4868 4217 4924
rect 4217 4868 4221 4924
rect 4157 4864 4221 4868
rect 9848 4924 9912 4928
rect 9848 4868 9852 4924
rect 9852 4868 9908 4924
rect 9908 4868 9912 4924
rect 9848 4864 9912 4868
rect 9928 4924 9992 4928
rect 9928 4868 9932 4924
rect 9932 4868 9988 4924
rect 9988 4868 9992 4924
rect 9928 4864 9992 4868
rect 10008 4924 10072 4928
rect 10008 4868 10012 4924
rect 10012 4868 10068 4924
rect 10068 4868 10072 4924
rect 10008 4864 10072 4868
rect 10088 4924 10152 4928
rect 10088 4868 10092 4924
rect 10092 4868 10148 4924
rect 10148 4868 10152 4924
rect 10088 4864 10152 4868
rect 15778 4924 15842 4928
rect 15778 4868 15782 4924
rect 15782 4868 15838 4924
rect 15838 4868 15842 4924
rect 15778 4864 15842 4868
rect 15858 4924 15922 4928
rect 15858 4868 15862 4924
rect 15862 4868 15918 4924
rect 15918 4868 15922 4924
rect 15858 4864 15922 4868
rect 15938 4924 16002 4928
rect 15938 4868 15942 4924
rect 15942 4868 15998 4924
rect 15998 4868 16002 4924
rect 15938 4864 16002 4868
rect 16018 4924 16082 4928
rect 16018 4868 16022 4924
rect 16022 4868 16078 4924
rect 16078 4868 16082 4924
rect 16018 4864 16082 4868
rect 6882 4380 6946 4384
rect 6882 4324 6886 4380
rect 6886 4324 6942 4380
rect 6942 4324 6946 4380
rect 6882 4320 6946 4324
rect 6962 4380 7026 4384
rect 6962 4324 6966 4380
rect 6966 4324 7022 4380
rect 7022 4324 7026 4380
rect 6962 4320 7026 4324
rect 7042 4380 7106 4384
rect 7042 4324 7046 4380
rect 7046 4324 7102 4380
rect 7102 4324 7106 4380
rect 7042 4320 7106 4324
rect 7122 4380 7186 4384
rect 7122 4324 7126 4380
rect 7126 4324 7182 4380
rect 7182 4324 7186 4380
rect 7122 4320 7186 4324
rect 12813 4380 12877 4384
rect 12813 4324 12817 4380
rect 12817 4324 12873 4380
rect 12873 4324 12877 4380
rect 12813 4320 12877 4324
rect 12893 4380 12957 4384
rect 12893 4324 12897 4380
rect 12897 4324 12953 4380
rect 12953 4324 12957 4380
rect 12893 4320 12957 4324
rect 12973 4380 13037 4384
rect 12973 4324 12977 4380
rect 12977 4324 13033 4380
rect 13033 4324 13037 4380
rect 12973 4320 13037 4324
rect 13053 4380 13117 4384
rect 13053 4324 13057 4380
rect 13057 4324 13113 4380
rect 13113 4324 13117 4380
rect 13053 4320 13117 4324
rect 3917 3836 3981 3840
rect 3917 3780 3921 3836
rect 3921 3780 3977 3836
rect 3977 3780 3981 3836
rect 3917 3776 3981 3780
rect 3997 3836 4061 3840
rect 3997 3780 4001 3836
rect 4001 3780 4057 3836
rect 4057 3780 4061 3836
rect 3997 3776 4061 3780
rect 4077 3836 4141 3840
rect 4077 3780 4081 3836
rect 4081 3780 4137 3836
rect 4137 3780 4141 3836
rect 4077 3776 4141 3780
rect 4157 3836 4221 3840
rect 4157 3780 4161 3836
rect 4161 3780 4217 3836
rect 4217 3780 4221 3836
rect 4157 3776 4221 3780
rect 9848 3836 9912 3840
rect 9848 3780 9852 3836
rect 9852 3780 9908 3836
rect 9908 3780 9912 3836
rect 9848 3776 9912 3780
rect 9928 3836 9992 3840
rect 9928 3780 9932 3836
rect 9932 3780 9988 3836
rect 9988 3780 9992 3836
rect 9928 3776 9992 3780
rect 10008 3836 10072 3840
rect 10008 3780 10012 3836
rect 10012 3780 10068 3836
rect 10068 3780 10072 3836
rect 10008 3776 10072 3780
rect 10088 3836 10152 3840
rect 10088 3780 10092 3836
rect 10092 3780 10148 3836
rect 10148 3780 10152 3836
rect 10088 3776 10152 3780
rect 15778 3836 15842 3840
rect 15778 3780 15782 3836
rect 15782 3780 15838 3836
rect 15838 3780 15842 3836
rect 15778 3776 15842 3780
rect 15858 3836 15922 3840
rect 15858 3780 15862 3836
rect 15862 3780 15918 3836
rect 15918 3780 15922 3836
rect 15858 3776 15922 3780
rect 15938 3836 16002 3840
rect 15938 3780 15942 3836
rect 15942 3780 15998 3836
rect 15998 3780 16002 3836
rect 15938 3776 16002 3780
rect 16018 3836 16082 3840
rect 16018 3780 16022 3836
rect 16022 3780 16078 3836
rect 16078 3780 16082 3836
rect 16018 3776 16082 3780
rect 6882 3292 6946 3296
rect 6882 3236 6886 3292
rect 6886 3236 6942 3292
rect 6942 3236 6946 3292
rect 6882 3232 6946 3236
rect 6962 3292 7026 3296
rect 6962 3236 6966 3292
rect 6966 3236 7022 3292
rect 7022 3236 7026 3292
rect 6962 3232 7026 3236
rect 7042 3292 7106 3296
rect 7042 3236 7046 3292
rect 7046 3236 7102 3292
rect 7102 3236 7106 3292
rect 7042 3232 7106 3236
rect 7122 3292 7186 3296
rect 7122 3236 7126 3292
rect 7126 3236 7182 3292
rect 7182 3236 7186 3292
rect 7122 3232 7186 3236
rect 12813 3292 12877 3296
rect 12813 3236 12817 3292
rect 12817 3236 12873 3292
rect 12873 3236 12877 3292
rect 12813 3232 12877 3236
rect 12893 3292 12957 3296
rect 12893 3236 12897 3292
rect 12897 3236 12953 3292
rect 12953 3236 12957 3292
rect 12893 3232 12957 3236
rect 12973 3292 13037 3296
rect 12973 3236 12977 3292
rect 12977 3236 13033 3292
rect 13033 3236 13037 3292
rect 12973 3232 13037 3236
rect 13053 3292 13117 3296
rect 13053 3236 13057 3292
rect 13057 3236 13113 3292
rect 13113 3236 13117 3292
rect 13053 3232 13117 3236
rect 16620 2892 16684 2956
rect 3917 2748 3981 2752
rect 3917 2692 3921 2748
rect 3921 2692 3977 2748
rect 3977 2692 3981 2748
rect 3917 2688 3981 2692
rect 3997 2748 4061 2752
rect 3997 2692 4001 2748
rect 4001 2692 4057 2748
rect 4057 2692 4061 2748
rect 3997 2688 4061 2692
rect 4077 2748 4141 2752
rect 4077 2692 4081 2748
rect 4081 2692 4137 2748
rect 4137 2692 4141 2748
rect 4077 2688 4141 2692
rect 4157 2748 4221 2752
rect 4157 2692 4161 2748
rect 4161 2692 4217 2748
rect 4217 2692 4221 2748
rect 4157 2688 4221 2692
rect 9848 2748 9912 2752
rect 9848 2692 9852 2748
rect 9852 2692 9908 2748
rect 9908 2692 9912 2748
rect 9848 2688 9912 2692
rect 9928 2748 9992 2752
rect 9928 2692 9932 2748
rect 9932 2692 9988 2748
rect 9988 2692 9992 2748
rect 9928 2688 9992 2692
rect 10008 2748 10072 2752
rect 10008 2692 10012 2748
rect 10012 2692 10068 2748
rect 10068 2692 10072 2748
rect 10008 2688 10072 2692
rect 10088 2748 10152 2752
rect 10088 2692 10092 2748
rect 10092 2692 10148 2748
rect 10148 2692 10152 2748
rect 10088 2688 10152 2692
rect 15778 2748 15842 2752
rect 15778 2692 15782 2748
rect 15782 2692 15838 2748
rect 15838 2692 15842 2748
rect 15778 2688 15842 2692
rect 15858 2748 15922 2752
rect 15858 2692 15862 2748
rect 15862 2692 15918 2748
rect 15918 2692 15922 2748
rect 15858 2688 15922 2692
rect 15938 2748 16002 2752
rect 15938 2692 15942 2748
rect 15942 2692 15998 2748
rect 15998 2692 16002 2748
rect 15938 2688 16002 2692
rect 16018 2748 16082 2752
rect 16018 2692 16022 2748
rect 16022 2692 16078 2748
rect 16078 2692 16082 2748
rect 16018 2688 16082 2692
rect 6882 2204 6946 2208
rect 6882 2148 6886 2204
rect 6886 2148 6942 2204
rect 6942 2148 6946 2204
rect 6882 2144 6946 2148
rect 6962 2204 7026 2208
rect 6962 2148 6966 2204
rect 6966 2148 7022 2204
rect 7022 2148 7026 2204
rect 6962 2144 7026 2148
rect 7042 2204 7106 2208
rect 7042 2148 7046 2204
rect 7046 2148 7102 2204
rect 7102 2148 7106 2204
rect 7042 2144 7106 2148
rect 7122 2204 7186 2208
rect 7122 2148 7126 2204
rect 7126 2148 7182 2204
rect 7182 2148 7186 2204
rect 7122 2144 7186 2148
rect 12813 2204 12877 2208
rect 12813 2148 12817 2204
rect 12817 2148 12873 2204
rect 12873 2148 12877 2204
rect 12813 2144 12877 2148
rect 12893 2204 12957 2208
rect 12893 2148 12897 2204
rect 12897 2148 12953 2204
rect 12953 2148 12957 2204
rect 12893 2144 12957 2148
rect 12973 2204 13037 2208
rect 12973 2148 12977 2204
rect 12977 2148 13033 2204
rect 13033 2148 13037 2204
rect 12973 2144 13037 2148
rect 13053 2204 13117 2208
rect 13053 2148 13057 2204
rect 13057 2148 13113 2204
rect 13113 2148 13117 2204
rect 13053 2144 13117 2148
<< metal4 >>
rect 3909 47360 4230 47376
rect 3909 47296 3917 47360
rect 3981 47296 3997 47360
rect 4061 47296 4077 47360
rect 4141 47296 4157 47360
rect 4221 47296 4230 47360
rect 3909 46272 4230 47296
rect 3909 46208 3917 46272
rect 3981 46208 3997 46272
rect 4061 46208 4077 46272
rect 4141 46208 4157 46272
rect 4221 46208 4230 46272
rect 3909 45184 4230 46208
rect 3909 45120 3917 45184
rect 3981 45120 3997 45184
rect 4061 45120 4077 45184
rect 4141 45120 4157 45184
rect 4221 45120 4230 45184
rect 3909 44096 4230 45120
rect 3909 44032 3917 44096
rect 3981 44032 3997 44096
rect 4061 44032 4077 44096
rect 4141 44032 4157 44096
rect 4221 44032 4230 44096
rect 3909 43008 4230 44032
rect 3909 42944 3917 43008
rect 3981 42944 3997 43008
rect 4061 42944 4077 43008
rect 4141 42944 4157 43008
rect 4221 42944 4230 43008
rect 3909 41920 4230 42944
rect 3909 41856 3917 41920
rect 3981 41856 3997 41920
rect 4061 41856 4077 41920
rect 4141 41856 4157 41920
rect 4221 41856 4230 41920
rect 3909 40832 4230 41856
rect 3909 40768 3917 40832
rect 3981 40768 3997 40832
rect 4061 40768 4077 40832
rect 4141 40768 4157 40832
rect 4221 40768 4230 40832
rect 3909 39744 4230 40768
rect 3909 39680 3917 39744
rect 3981 39680 3997 39744
rect 4061 39680 4077 39744
rect 4141 39680 4157 39744
rect 4221 39680 4230 39744
rect 3909 38656 4230 39680
rect 3909 38592 3917 38656
rect 3981 38592 3997 38656
rect 4061 38592 4077 38656
rect 4141 38592 4157 38656
rect 4221 38592 4230 38656
rect 3909 37568 4230 38592
rect 3909 37504 3917 37568
rect 3981 37504 3997 37568
rect 4061 37504 4077 37568
rect 4141 37504 4157 37568
rect 4221 37504 4230 37568
rect 3909 36480 4230 37504
rect 3909 36416 3917 36480
rect 3981 36416 3997 36480
rect 4061 36416 4077 36480
rect 4141 36416 4157 36480
rect 4221 36416 4230 36480
rect 3909 35392 4230 36416
rect 3909 35328 3917 35392
rect 3981 35328 3997 35392
rect 4061 35328 4077 35392
rect 4141 35328 4157 35392
rect 4221 35328 4230 35392
rect 3909 34304 4230 35328
rect 3909 34240 3917 34304
rect 3981 34240 3997 34304
rect 4061 34240 4077 34304
rect 4141 34240 4157 34304
rect 4221 34240 4230 34304
rect 3909 33216 4230 34240
rect 3909 33152 3917 33216
rect 3981 33152 3997 33216
rect 4061 33152 4077 33216
rect 4141 33152 4157 33216
rect 4221 33152 4230 33216
rect 3909 32128 4230 33152
rect 3909 32064 3917 32128
rect 3981 32064 3997 32128
rect 4061 32064 4077 32128
rect 4141 32064 4157 32128
rect 4221 32064 4230 32128
rect 3909 31040 4230 32064
rect 3909 30976 3917 31040
rect 3981 30976 3997 31040
rect 4061 30976 4077 31040
rect 4141 30976 4157 31040
rect 4221 30976 4230 31040
rect 3909 29952 4230 30976
rect 3909 29888 3917 29952
rect 3981 29888 3997 29952
rect 4061 29888 4077 29952
rect 4141 29888 4157 29952
rect 4221 29888 4230 29952
rect 3909 28864 4230 29888
rect 3909 28800 3917 28864
rect 3981 28800 3997 28864
rect 4061 28800 4077 28864
rect 4141 28800 4157 28864
rect 4221 28800 4230 28864
rect 3909 27776 4230 28800
rect 3909 27712 3917 27776
rect 3981 27712 3997 27776
rect 4061 27712 4077 27776
rect 4141 27712 4157 27776
rect 4221 27712 4230 27776
rect 3909 26688 4230 27712
rect 3909 26624 3917 26688
rect 3981 26624 3997 26688
rect 4061 26624 4077 26688
rect 4141 26624 4157 26688
rect 4221 26624 4230 26688
rect 3909 25600 4230 26624
rect 3909 25536 3917 25600
rect 3981 25536 3997 25600
rect 4061 25536 4077 25600
rect 4141 25536 4157 25600
rect 4221 25536 4230 25600
rect 3909 24512 4230 25536
rect 3909 24448 3917 24512
rect 3981 24448 3997 24512
rect 4061 24448 4077 24512
rect 4141 24448 4157 24512
rect 4221 24448 4230 24512
rect 3909 23424 4230 24448
rect 3909 23360 3917 23424
rect 3981 23360 3997 23424
rect 4061 23360 4077 23424
rect 4141 23360 4157 23424
rect 4221 23360 4230 23424
rect 3909 22336 4230 23360
rect 3909 22272 3917 22336
rect 3981 22272 3997 22336
rect 4061 22272 4077 22336
rect 4141 22272 4157 22336
rect 4221 22272 4230 22336
rect 3909 21248 4230 22272
rect 3909 21184 3917 21248
rect 3981 21184 3997 21248
rect 4061 21184 4077 21248
rect 4141 21184 4157 21248
rect 4221 21184 4230 21248
rect 3909 20160 4230 21184
rect 3909 20096 3917 20160
rect 3981 20096 3997 20160
rect 4061 20096 4077 20160
rect 4141 20096 4157 20160
rect 4221 20096 4230 20160
rect 3909 19072 4230 20096
rect 3909 19008 3917 19072
rect 3981 19008 3997 19072
rect 4061 19008 4077 19072
rect 4141 19008 4157 19072
rect 4221 19008 4230 19072
rect 3909 17984 4230 19008
rect 3909 17920 3917 17984
rect 3981 17920 3997 17984
rect 4061 17920 4077 17984
rect 4141 17920 4157 17984
rect 4221 17920 4230 17984
rect 3909 16896 4230 17920
rect 3909 16832 3917 16896
rect 3981 16832 3997 16896
rect 4061 16832 4077 16896
rect 4141 16832 4157 16896
rect 4221 16832 4230 16896
rect 3909 15808 4230 16832
rect 3909 15744 3917 15808
rect 3981 15744 3997 15808
rect 4061 15744 4077 15808
rect 4141 15744 4157 15808
rect 4221 15744 4230 15808
rect 3909 14720 4230 15744
rect 3909 14656 3917 14720
rect 3981 14656 3997 14720
rect 4061 14656 4077 14720
rect 4141 14656 4157 14720
rect 4221 14656 4230 14720
rect 3909 13632 4230 14656
rect 3909 13568 3917 13632
rect 3981 13568 3997 13632
rect 4061 13568 4077 13632
rect 4141 13568 4157 13632
rect 4221 13568 4230 13632
rect 3909 12544 4230 13568
rect 3909 12480 3917 12544
rect 3981 12480 3997 12544
rect 4061 12480 4077 12544
rect 4141 12480 4157 12544
rect 4221 12480 4230 12544
rect 3909 11456 4230 12480
rect 3909 11392 3917 11456
rect 3981 11392 3997 11456
rect 4061 11392 4077 11456
rect 4141 11392 4157 11456
rect 4221 11392 4230 11456
rect 3909 10368 4230 11392
rect 3909 10304 3917 10368
rect 3981 10304 3997 10368
rect 4061 10304 4077 10368
rect 4141 10304 4157 10368
rect 4221 10304 4230 10368
rect 3909 9280 4230 10304
rect 3909 9216 3917 9280
rect 3981 9216 3997 9280
rect 4061 9216 4077 9280
rect 4141 9216 4157 9280
rect 4221 9216 4230 9280
rect 3909 8192 4230 9216
rect 3909 8128 3917 8192
rect 3981 8128 3997 8192
rect 4061 8128 4077 8192
rect 4141 8128 4157 8192
rect 4221 8128 4230 8192
rect 3909 7104 4230 8128
rect 3909 7040 3917 7104
rect 3981 7040 3997 7104
rect 4061 7040 4077 7104
rect 4141 7040 4157 7104
rect 4221 7040 4230 7104
rect 3909 6016 4230 7040
rect 3909 5952 3917 6016
rect 3981 5952 3997 6016
rect 4061 5952 4077 6016
rect 4141 5952 4157 6016
rect 4221 5952 4230 6016
rect 3909 4928 4230 5952
rect 3909 4864 3917 4928
rect 3981 4864 3997 4928
rect 4061 4864 4077 4928
rect 4141 4864 4157 4928
rect 4221 4864 4230 4928
rect 3909 3840 4230 4864
rect 3909 3776 3917 3840
rect 3981 3776 3997 3840
rect 4061 3776 4077 3840
rect 4141 3776 4157 3840
rect 4221 3776 4230 3840
rect 3909 2752 4230 3776
rect 3909 2688 3917 2752
rect 3981 2688 3997 2752
rect 4061 2688 4077 2752
rect 4141 2688 4157 2752
rect 4221 2688 4230 2752
rect 3909 2128 4230 2688
rect 6874 46816 7194 47376
rect 6874 46752 6882 46816
rect 6946 46752 6962 46816
rect 7026 46752 7042 46816
rect 7106 46752 7122 46816
rect 7186 46752 7194 46816
rect 6874 45728 7194 46752
rect 6874 45664 6882 45728
rect 6946 45664 6962 45728
rect 7026 45664 7042 45728
rect 7106 45664 7122 45728
rect 7186 45664 7194 45728
rect 6874 44640 7194 45664
rect 6874 44576 6882 44640
rect 6946 44576 6962 44640
rect 7026 44576 7042 44640
rect 7106 44576 7122 44640
rect 7186 44576 7194 44640
rect 6874 43552 7194 44576
rect 6874 43488 6882 43552
rect 6946 43488 6962 43552
rect 7026 43488 7042 43552
rect 7106 43488 7122 43552
rect 7186 43488 7194 43552
rect 6874 42464 7194 43488
rect 6874 42400 6882 42464
rect 6946 42400 6962 42464
rect 7026 42400 7042 42464
rect 7106 42400 7122 42464
rect 7186 42400 7194 42464
rect 6874 41376 7194 42400
rect 6874 41312 6882 41376
rect 6946 41312 6962 41376
rect 7026 41312 7042 41376
rect 7106 41312 7122 41376
rect 7186 41312 7194 41376
rect 6874 40288 7194 41312
rect 6874 40224 6882 40288
rect 6946 40224 6962 40288
rect 7026 40224 7042 40288
rect 7106 40224 7122 40288
rect 7186 40224 7194 40288
rect 6874 39200 7194 40224
rect 6874 39136 6882 39200
rect 6946 39136 6962 39200
rect 7026 39136 7042 39200
rect 7106 39136 7122 39200
rect 7186 39136 7194 39200
rect 6874 38112 7194 39136
rect 6874 38048 6882 38112
rect 6946 38048 6962 38112
rect 7026 38048 7042 38112
rect 7106 38048 7122 38112
rect 7186 38048 7194 38112
rect 6874 37024 7194 38048
rect 6874 36960 6882 37024
rect 6946 36960 6962 37024
rect 7026 36960 7042 37024
rect 7106 36960 7122 37024
rect 7186 36960 7194 37024
rect 6874 35936 7194 36960
rect 6874 35872 6882 35936
rect 6946 35872 6962 35936
rect 7026 35872 7042 35936
rect 7106 35872 7122 35936
rect 7186 35872 7194 35936
rect 6874 34848 7194 35872
rect 6874 34784 6882 34848
rect 6946 34784 6962 34848
rect 7026 34784 7042 34848
rect 7106 34784 7122 34848
rect 7186 34784 7194 34848
rect 6874 33760 7194 34784
rect 6874 33696 6882 33760
rect 6946 33696 6962 33760
rect 7026 33696 7042 33760
rect 7106 33696 7122 33760
rect 7186 33696 7194 33760
rect 6874 32672 7194 33696
rect 6874 32608 6882 32672
rect 6946 32608 6962 32672
rect 7026 32608 7042 32672
rect 7106 32608 7122 32672
rect 7186 32608 7194 32672
rect 6874 31584 7194 32608
rect 6874 31520 6882 31584
rect 6946 31520 6962 31584
rect 7026 31520 7042 31584
rect 7106 31520 7122 31584
rect 7186 31520 7194 31584
rect 6874 30496 7194 31520
rect 6874 30432 6882 30496
rect 6946 30432 6962 30496
rect 7026 30432 7042 30496
rect 7106 30432 7122 30496
rect 7186 30432 7194 30496
rect 6874 29408 7194 30432
rect 6874 29344 6882 29408
rect 6946 29344 6962 29408
rect 7026 29344 7042 29408
rect 7106 29344 7122 29408
rect 7186 29344 7194 29408
rect 6874 28320 7194 29344
rect 6874 28256 6882 28320
rect 6946 28256 6962 28320
rect 7026 28256 7042 28320
rect 7106 28256 7122 28320
rect 7186 28256 7194 28320
rect 6874 27232 7194 28256
rect 6874 27168 6882 27232
rect 6946 27168 6962 27232
rect 7026 27168 7042 27232
rect 7106 27168 7122 27232
rect 7186 27168 7194 27232
rect 6874 26144 7194 27168
rect 6874 26080 6882 26144
rect 6946 26080 6962 26144
rect 7026 26080 7042 26144
rect 7106 26080 7122 26144
rect 7186 26080 7194 26144
rect 6874 25056 7194 26080
rect 6874 24992 6882 25056
rect 6946 24992 6962 25056
rect 7026 24992 7042 25056
rect 7106 24992 7122 25056
rect 7186 24992 7194 25056
rect 6874 23968 7194 24992
rect 6874 23904 6882 23968
rect 6946 23904 6962 23968
rect 7026 23904 7042 23968
rect 7106 23904 7122 23968
rect 7186 23904 7194 23968
rect 6874 22880 7194 23904
rect 6874 22816 6882 22880
rect 6946 22816 6962 22880
rect 7026 22816 7042 22880
rect 7106 22816 7122 22880
rect 7186 22816 7194 22880
rect 6874 21792 7194 22816
rect 6874 21728 6882 21792
rect 6946 21728 6962 21792
rect 7026 21728 7042 21792
rect 7106 21728 7122 21792
rect 7186 21728 7194 21792
rect 6874 20704 7194 21728
rect 6874 20640 6882 20704
rect 6946 20640 6962 20704
rect 7026 20640 7042 20704
rect 7106 20640 7122 20704
rect 7186 20640 7194 20704
rect 6874 19616 7194 20640
rect 6874 19552 6882 19616
rect 6946 19552 6962 19616
rect 7026 19552 7042 19616
rect 7106 19552 7122 19616
rect 7186 19552 7194 19616
rect 6874 18528 7194 19552
rect 6874 18464 6882 18528
rect 6946 18464 6962 18528
rect 7026 18464 7042 18528
rect 7106 18464 7122 18528
rect 7186 18464 7194 18528
rect 6874 17440 7194 18464
rect 6874 17376 6882 17440
rect 6946 17376 6962 17440
rect 7026 17376 7042 17440
rect 7106 17376 7122 17440
rect 7186 17376 7194 17440
rect 6874 16352 7194 17376
rect 6874 16288 6882 16352
rect 6946 16288 6962 16352
rect 7026 16288 7042 16352
rect 7106 16288 7122 16352
rect 7186 16288 7194 16352
rect 6874 15264 7194 16288
rect 6874 15200 6882 15264
rect 6946 15200 6962 15264
rect 7026 15200 7042 15264
rect 7106 15200 7122 15264
rect 7186 15200 7194 15264
rect 6874 14176 7194 15200
rect 6874 14112 6882 14176
rect 6946 14112 6962 14176
rect 7026 14112 7042 14176
rect 7106 14112 7122 14176
rect 7186 14112 7194 14176
rect 6874 13088 7194 14112
rect 6874 13024 6882 13088
rect 6946 13024 6962 13088
rect 7026 13024 7042 13088
rect 7106 13024 7122 13088
rect 7186 13024 7194 13088
rect 6874 12000 7194 13024
rect 6874 11936 6882 12000
rect 6946 11936 6962 12000
rect 7026 11936 7042 12000
rect 7106 11936 7122 12000
rect 7186 11936 7194 12000
rect 6874 10912 7194 11936
rect 6874 10848 6882 10912
rect 6946 10848 6962 10912
rect 7026 10848 7042 10912
rect 7106 10848 7122 10912
rect 7186 10848 7194 10912
rect 6874 9824 7194 10848
rect 6874 9760 6882 9824
rect 6946 9760 6962 9824
rect 7026 9760 7042 9824
rect 7106 9760 7122 9824
rect 7186 9760 7194 9824
rect 6874 8736 7194 9760
rect 6874 8672 6882 8736
rect 6946 8672 6962 8736
rect 7026 8672 7042 8736
rect 7106 8672 7122 8736
rect 7186 8672 7194 8736
rect 6874 7648 7194 8672
rect 6874 7584 6882 7648
rect 6946 7584 6962 7648
rect 7026 7584 7042 7648
rect 7106 7584 7122 7648
rect 7186 7584 7194 7648
rect 6874 6560 7194 7584
rect 6874 6496 6882 6560
rect 6946 6496 6962 6560
rect 7026 6496 7042 6560
rect 7106 6496 7122 6560
rect 7186 6496 7194 6560
rect 6874 5472 7194 6496
rect 6874 5408 6882 5472
rect 6946 5408 6962 5472
rect 7026 5408 7042 5472
rect 7106 5408 7122 5472
rect 7186 5408 7194 5472
rect 6874 4384 7194 5408
rect 6874 4320 6882 4384
rect 6946 4320 6962 4384
rect 7026 4320 7042 4384
rect 7106 4320 7122 4384
rect 7186 4320 7194 4384
rect 6874 3296 7194 4320
rect 6874 3232 6882 3296
rect 6946 3232 6962 3296
rect 7026 3232 7042 3296
rect 7106 3232 7122 3296
rect 7186 3232 7194 3296
rect 6874 2208 7194 3232
rect 6874 2144 6882 2208
rect 6946 2144 6962 2208
rect 7026 2144 7042 2208
rect 7106 2144 7122 2208
rect 7186 2144 7194 2208
rect 6874 2128 7194 2144
rect 9840 47360 10160 47376
rect 9840 47296 9848 47360
rect 9912 47296 9928 47360
rect 9992 47296 10008 47360
rect 10072 47296 10088 47360
rect 10152 47296 10160 47360
rect 9840 46272 10160 47296
rect 9840 46208 9848 46272
rect 9912 46208 9928 46272
rect 9992 46208 10008 46272
rect 10072 46208 10088 46272
rect 10152 46208 10160 46272
rect 9840 45184 10160 46208
rect 9840 45120 9848 45184
rect 9912 45120 9928 45184
rect 9992 45120 10008 45184
rect 10072 45120 10088 45184
rect 10152 45120 10160 45184
rect 9840 44096 10160 45120
rect 9840 44032 9848 44096
rect 9912 44032 9928 44096
rect 9992 44032 10008 44096
rect 10072 44032 10088 44096
rect 10152 44032 10160 44096
rect 9840 43008 10160 44032
rect 9840 42944 9848 43008
rect 9912 42944 9928 43008
rect 9992 42944 10008 43008
rect 10072 42944 10088 43008
rect 10152 42944 10160 43008
rect 9840 41920 10160 42944
rect 9840 41856 9848 41920
rect 9912 41856 9928 41920
rect 9992 41856 10008 41920
rect 10072 41856 10088 41920
rect 10152 41856 10160 41920
rect 9840 40832 10160 41856
rect 9840 40768 9848 40832
rect 9912 40768 9928 40832
rect 9992 40768 10008 40832
rect 10072 40768 10088 40832
rect 10152 40768 10160 40832
rect 9840 39744 10160 40768
rect 9840 39680 9848 39744
rect 9912 39680 9928 39744
rect 9992 39680 10008 39744
rect 10072 39680 10088 39744
rect 10152 39680 10160 39744
rect 9840 38656 10160 39680
rect 9840 38592 9848 38656
rect 9912 38592 9928 38656
rect 9992 38592 10008 38656
rect 10072 38592 10088 38656
rect 10152 38592 10160 38656
rect 9840 37568 10160 38592
rect 9840 37504 9848 37568
rect 9912 37504 9928 37568
rect 9992 37504 10008 37568
rect 10072 37504 10088 37568
rect 10152 37504 10160 37568
rect 9840 36480 10160 37504
rect 9840 36416 9848 36480
rect 9912 36416 9928 36480
rect 9992 36416 10008 36480
rect 10072 36416 10088 36480
rect 10152 36416 10160 36480
rect 9840 35392 10160 36416
rect 9840 35328 9848 35392
rect 9912 35328 9928 35392
rect 9992 35328 10008 35392
rect 10072 35328 10088 35392
rect 10152 35328 10160 35392
rect 9840 34304 10160 35328
rect 9840 34240 9848 34304
rect 9912 34240 9928 34304
rect 9992 34240 10008 34304
rect 10072 34240 10088 34304
rect 10152 34240 10160 34304
rect 9840 33216 10160 34240
rect 9840 33152 9848 33216
rect 9912 33152 9928 33216
rect 9992 33152 10008 33216
rect 10072 33152 10088 33216
rect 10152 33152 10160 33216
rect 9840 32128 10160 33152
rect 9840 32064 9848 32128
rect 9912 32064 9928 32128
rect 9992 32064 10008 32128
rect 10072 32064 10088 32128
rect 10152 32064 10160 32128
rect 9840 31040 10160 32064
rect 9840 30976 9848 31040
rect 9912 30976 9928 31040
rect 9992 30976 10008 31040
rect 10072 30976 10088 31040
rect 10152 30976 10160 31040
rect 9840 29952 10160 30976
rect 9840 29888 9848 29952
rect 9912 29888 9928 29952
rect 9992 29888 10008 29952
rect 10072 29888 10088 29952
rect 10152 29888 10160 29952
rect 9840 28864 10160 29888
rect 9840 28800 9848 28864
rect 9912 28800 9928 28864
rect 9992 28800 10008 28864
rect 10072 28800 10088 28864
rect 10152 28800 10160 28864
rect 9840 27776 10160 28800
rect 9840 27712 9848 27776
rect 9912 27712 9928 27776
rect 9992 27712 10008 27776
rect 10072 27712 10088 27776
rect 10152 27712 10160 27776
rect 9840 26688 10160 27712
rect 9840 26624 9848 26688
rect 9912 26624 9928 26688
rect 9992 26624 10008 26688
rect 10072 26624 10088 26688
rect 10152 26624 10160 26688
rect 9840 25600 10160 26624
rect 9840 25536 9848 25600
rect 9912 25536 9928 25600
rect 9992 25536 10008 25600
rect 10072 25536 10088 25600
rect 10152 25536 10160 25600
rect 9840 24512 10160 25536
rect 9840 24448 9848 24512
rect 9912 24448 9928 24512
rect 9992 24448 10008 24512
rect 10072 24448 10088 24512
rect 10152 24448 10160 24512
rect 9840 23424 10160 24448
rect 9840 23360 9848 23424
rect 9912 23360 9928 23424
rect 9992 23360 10008 23424
rect 10072 23360 10088 23424
rect 10152 23360 10160 23424
rect 9840 22336 10160 23360
rect 9840 22272 9848 22336
rect 9912 22272 9928 22336
rect 9992 22272 10008 22336
rect 10072 22272 10088 22336
rect 10152 22272 10160 22336
rect 9840 21248 10160 22272
rect 9840 21184 9848 21248
rect 9912 21184 9928 21248
rect 9992 21184 10008 21248
rect 10072 21184 10088 21248
rect 10152 21184 10160 21248
rect 9840 20160 10160 21184
rect 9840 20096 9848 20160
rect 9912 20096 9928 20160
rect 9992 20096 10008 20160
rect 10072 20096 10088 20160
rect 10152 20096 10160 20160
rect 9840 19072 10160 20096
rect 9840 19008 9848 19072
rect 9912 19008 9928 19072
rect 9992 19008 10008 19072
rect 10072 19008 10088 19072
rect 10152 19008 10160 19072
rect 9840 17984 10160 19008
rect 9840 17920 9848 17984
rect 9912 17920 9928 17984
rect 9992 17920 10008 17984
rect 10072 17920 10088 17984
rect 10152 17920 10160 17984
rect 9840 16896 10160 17920
rect 9840 16832 9848 16896
rect 9912 16832 9928 16896
rect 9992 16832 10008 16896
rect 10072 16832 10088 16896
rect 10152 16832 10160 16896
rect 9840 15808 10160 16832
rect 9840 15744 9848 15808
rect 9912 15744 9928 15808
rect 9992 15744 10008 15808
rect 10072 15744 10088 15808
rect 10152 15744 10160 15808
rect 9840 14720 10160 15744
rect 9840 14656 9848 14720
rect 9912 14656 9928 14720
rect 9992 14656 10008 14720
rect 10072 14656 10088 14720
rect 10152 14656 10160 14720
rect 9840 13632 10160 14656
rect 9840 13568 9848 13632
rect 9912 13568 9928 13632
rect 9992 13568 10008 13632
rect 10072 13568 10088 13632
rect 10152 13568 10160 13632
rect 9840 12544 10160 13568
rect 9840 12480 9848 12544
rect 9912 12480 9928 12544
rect 9992 12480 10008 12544
rect 10072 12480 10088 12544
rect 10152 12480 10160 12544
rect 9840 11456 10160 12480
rect 9840 11392 9848 11456
rect 9912 11392 9928 11456
rect 9992 11392 10008 11456
rect 10072 11392 10088 11456
rect 10152 11392 10160 11456
rect 9840 10368 10160 11392
rect 9840 10304 9848 10368
rect 9912 10304 9928 10368
rect 9992 10304 10008 10368
rect 10072 10304 10088 10368
rect 10152 10304 10160 10368
rect 9840 9280 10160 10304
rect 9840 9216 9848 9280
rect 9912 9216 9928 9280
rect 9992 9216 10008 9280
rect 10072 9216 10088 9280
rect 10152 9216 10160 9280
rect 9840 8192 10160 9216
rect 9840 8128 9848 8192
rect 9912 8128 9928 8192
rect 9992 8128 10008 8192
rect 10072 8128 10088 8192
rect 10152 8128 10160 8192
rect 9840 7104 10160 8128
rect 9840 7040 9848 7104
rect 9912 7040 9928 7104
rect 9992 7040 10008 7104
rect 10072 7040 10088 7104
rect 10152 7040 10160 7104
rect 9840 6016 10160 7040
rect 9840 5952 9848 6016
rect 9912 5952 9928 6016
rect 9992 5952 10008 6016
rect 10072 5952 10088 6016
rect 10152 5952 10160 6016
rect 9840 4928 10160 5952
rect 9840 4864 9848 4928
rect 9912 4864 9928 4928
rect 9992 4864 10008 4928
rect 10072 4864 10088 4928
rect 10152 4864 10160 4928
rect 9840 3840 10160 4864
rect 9840 3776 9848 3840
rect 9912 3776 9928 3840
rect 9992 3776 10008 3840
rect 10072 3776 10088 3840
rect 10152 3776 10160 3840
rect 9840 2752 10160 3776
rect 9840 2688 9848 2752
rect 9912 2688 9928 2752
rect 9992 2688 10008 2752
rect 10072 2688 10088 2752
rect 10152 2688 10160 2752
rect 9840 2128 10160 2688
rect 12805 46816 13125 47376
rect 12805 46752 12813 46816
rect 12877 46752 12893 46816
rect 12957 46752 12973 46816
rect 13037 46752 13053 46816
rect 13117 46752 13125 46816
rect 12805 45728 13125 46752
rect 15770 47360 16091 47376
rect 15770 47296 15778 47360
rect 15842 47296 15858 47360
rect 15922 47296 15938 47360
rect 16002 47296 16018 47360
rect 16082 47296 16091 47360
rect 15770 46272 16091 47296
rect 15770 46208 15778 46272
rect 15842 46208 15858 46272
rect 15922 46208 15938 46272
rect 16002 46208 16018 46272
rect 16082 46208 16091 46272
rect 15515 45932 15581 45933
rect 15515 45868 15516 45932
rect 15580 45868 15581 45932
rect 15515 45867 15581 45868
rect 12805 45664 12813 45728
rect 12877 45664 12893 45728
rect 12957 45664 12973 45728
rect 13037 45664 13053 45728
rect 13117 45664 13125 45728
rect 12805 44640 13125 45664
rect 12805 44576 12813 44640
rect 12877 44576 12893 44640
rect 12957 44576 12973 44640
rect 13037 44576 13053 44640
rect 13117 44576 13125 44640
rect 12805 43552 13125 44576
rect 12805 43488 12813 43552
rect 12877 43488 12893 43552
rect 12957 43488 12973 43552
rect 13037 43488 13053 43552
rect 13117 43488 13125 43552
rect 12805 42464 13125 43488
rect 12805 42400 12813 42464
rect 12877 42400 12893 42464
rect 12957 42400 12973 42464
rect 13037 42400 13053 42464
rect 13117 42400 13125 42464
rect 12805 41376 13125 42400
rect 12805 41312 12813 41376
rect 12877 41312 12893 41376
rect 12957 41312 12973 41376
rect 13037 41312 13053 41376
rect 13117 41312 13125 41376
rect 12805 40288 13125 41312
rect 12805 40224 12813 40288
rect 12877 40224 12893 40288
rect 12957 40224 12973 40288
rect 13037 40224 13053 40288
rect 13117 40224 13125 40288
rect 12805 39200 13125 40224
rect 12805 39136 12813 39200
rect 12877 39136 12893 39200
rect 12957 39136 12973 39200
rect 13037 39136 13053 39200
rect 13117 39136 13125 39200
rect 12805 38112 13125 39136
rect 12805 38048 12813 38112
rect 12877 38048 12893 38112
rect 12957 38048 12973 38112
rect 13037 38048 13053 38112
rect 13117 38048 13125 38112
rect 12805 37024 13125 38048
rect 12805 36960 12813 37024
rect 12877 36960 12893 37024
rect 12957 36960 12973 37024
rect 13037 36960 13053 37024
rect 13117 36960 13125 37024
rect 12805 35936 13125 36960
rect 12805 35872 12813 35936
rect 12877 35872 12893 35936
rect 12957 35872 12973 35936
rect 13037 35872 13053 35936
rect 13117 35872 13125 35936
rect 12805 34848 13125 35872
rect 12805 34784 12813 34848
rect 12877 34784 12893 34848
rect 12957 34784 12973 34848
rect 13037 34784 13053 34848
rect 13117 34784 13125 34848
rect 12805 33760 13125 34784
rect 12805 33696 12813 33760
rect 12877 33696 12893 33760
rect 12957 33696 12973 33760
rect 13037 33696 13053 33760
rect 13117 33696 13125 33760
rect 12805 32672 13125 33696
rect 12805 32608 12813 32672
rect 12877 32608 12893 32672
rect 12957 32608 12973 32672
rect 13037 32608 13053 32672
rect 13117 32608 13125 32672
rect 12805 31584 13125 32608
rect 12805 31520 12813 31584
rect 12877 31520 12893 31584
rect 12957 31520 12973 31584
rect 13037 31520 13053 31584
rect 13117 31520 13125 31584
rect 12805 30496 13125 31520
rect 12805 30432 12813 30496
rect 12877 30432 12893 30496
rect 12957 30432 12973 30496
rect 13037 30432 13053 30496
rect 13117 30432 13125 30496
rect 12805 29408 13125 30432
rect 12805 29344 12813 29408
rect 12877 29344 12893 29408
rect 12957 29344 12973 29408
rect 13037 29344 13053 29408
rect 13117 29344 13125 29408
rect 12805 28320 13125 29344
rect 12805 28256 12813 28320
rect 12877 28256 12893 28320
rect 12957 28256 12973 28320
rect 13037 28256 13053 28320
rect 13117 28256 13125 28320
rect 12805 27232 13125 28256
rect 12805 27168 12813 27232
rect 12877 27168 12893 27232
rect 12957 27168 12973 27232
rect 13037 27168 13053 27232
rect 13117 27168 13125 27232
rect 12805 26144 13125 27168
rect 12805 26080 12813 26144
rect 12877 26080 12893 26144
rect 12957 26080 12973 26144
rect 13037 26080 13053 26144
rect 13117 26080 13125 26144
rect 12805 25056 13125 26080
rect 15518 25533 15578 45867
rect 15770 45184 16091 46208
rect 15770 45120 15778 45184
rect 15842 45120 15858 45184
rect 15922 45120 15938 45184
rect 16002 45120 16018 45184
rect 16082 45120 16091 45184
rect 15770 44096 16091 45120
rect 15770 44032 15778 44096
rect 15842 44032 15858 44096
rect 15922 44032 15938 44096
rect 16002 44032 16018 44096
rect 16082 44032 16091 44096
rect 15770 43008 16091 44032
rect 15770 42944 15778 43008
rect 15842 42944 15858 43008
rect 15922 42944 15938 43008
rect 16002 42944 16018 43008
rect 16082 42944 16091 43008
rect 15770 41920 16091 42944
rect 15770 41856 15778 41920
rect 15842 41856 15858 41920
rect 15922 41856 15938 41920
rect 16002 41856 16018 41920
rect 16082 41856 16091 41920
rect 15770 40832 16091 41856
rect 15770 40768 15778 40832
rect 15842 40768 15858 40832
rect 15922 40768 15938 40832
rect 16002 40768 16018 40832
rect 16082 40768 16091 40832
rect 15770 39744 16091 40768
rect 15770 39680 15778 39744
rect 15842 39680 15858 39744
rect 15922 39680 15938 39744
rect 16002 39680 16018 39744
rect 16082 39680 16091 39744
rect 15770 38656 16091 39680
rect 15770 38592 15778 38656
rect 15842 38592 15858 38656
rect 15922 38592 15938 38656
rect 16002 38592 16018 38656
rect 16082 38592 16091 38656
rect 15770 37568 16091 38592
rect 15770 37504 15778 37568
rect 15842 37504 15858 37568
rect 15922 37504 15938 37568
rect 16002 37504 16018 37568
rect 16082 37504 16091 37568
rect 15770 36480 16091 37504
rect 15770 36416 15778 36480
rect 15842 36416 15858 36480
rect 15922 36416 15938 36480
rect 16002 36416 16018 36480
rect 16082 36416 16091 36480
rect 15770 35392 16091 36416
rect 15770 35328 15778 35392
rect 15842 35328 15858 35392
rect 15922 35328 15938 35392
rect 16002 35328 16018 35392
rect 16082 35328 16091 35392
rect 15770 34304 16091 35328
rect 15770 34240 15778 34304
rect 15842 34240 15858 34304
rect 15922 34240 15938 34304
rect 16002 34240 16018 34304
rect 16082 34240 16091 34304
rect 15770 33216 16091 34240
rect 16619 33284 16685 33285
rect 16619 33220 16620 33284
rect 16684 33220 16685 33284
rect 16619 33219 16685 33220
rect 15770 33152 15778 33216
rect 15842 33152 15858 33216
rect 15922 33152 15938 33216
rect 16002 33152 16018 33216
rect 16082 33152 16091 33216
rect 15770 32128 16091 33152
rect 15770 32064 15778 32128
rect 15842 32064 15858 32128
rect 15922 32064 15938 32128
rect 16002 32064 16018 32128
rect 16082 32064 16091 32128
rect 15770 31040 16091 32064
rect 15770 30976 15778 31040
rect 15842 30976 15858 31040
rect 15922 30976 15938 31040
rect 16002 30976 16018 31040
rect 16082 30976 16091 31040
rect 15770 29952 16091 30976
rect 15770 29888 15778 29952
rect 15842 29888 15858 29952
rect 15922 29888 15938 29952
rect 16002 29888 16018 29952
rect 16082 29888 16091 29952
rect 15770 28864 16091 29888
rect 15770 28800 15778 28864
rect 15842 28800 15858 28864
rect 15922 28800 15938 28864
rect 16002 28800 16018 28864
rect 16082 28800 16091 28864
rect 15770 27776 16091 28800
rect 15770 27712 15778 27776
rect 15842 27712 15858 27776
rect 15922 27712 15938 27776
rect 16002 27712 16018 27776
rect 16082 27712 16091 27776
rect 15770 26688 16091 27712
rect 15770 26624 15778 26688
rect 15842 26624 15858 26688
rect 15922 26624 15938 26688
rect 16002 26624 16018 26688
rect 16082 26624 16091 26688
rect 15770 25600 16091 26624
rect 15770 25536 15778 25600
rect 15842 25536 15858 25600
rect 15922 25536 15938 25600
rect 16002 25536 16018 25600
rect 16082 25536 16091 25600
rect 15515 25532 15581 25533
rect 15515 25468 15516 25532
rect 15580 25468 15581 25532
rect 15515 25467 15581 25468
rect 12805 24992 12813 25056
rect 12877 24992 12893 25056
rect 12957 24992 12973 25056
rect 13037 24992 13053 25056
rect 13117 24992 13125 25056
rect 12805 23968 13125 24992
rect 12805 23904 12813 23968
rect 12877 23904 12893 23968
rect 12957 23904 12973 23968
rect 13037 23904 13053 23968
rect 13117 23904 13125 23968
rect 12805 22880 13125 23904
rect 12805 22816 12813 22880
rect 12877 22816 12893 22880
rect 12957 22816 12973 22880
rect 13037 22816 13053 22880
rect 13117 22816 13125 22880
rect 12805 21792 13125 22816
rect 12805 21728 12813 21792
rect 12877 21728 12893 21792
rect 12957 21728 12973 21792
rect 13037 21728 13053 21792
rect 13117 21728 13125 21792
rect 12805 20704 13125 21728
rect 12805 20640 12813 20704
rect 12877 20640 12893 20704
rect 12957 20640 12973 20704
rect 13037 20640 13053 20704
rect 13117 20640 13125 20704
rect 12805 19616 13125 20640
rect 12805 19552 12813 19616
rect 12877 19552 12893 19616
rect 12957 19552 12973 19616
rect 13037 19552 13053 19616
rect 13117 19552 13125 19616
rect 12805 18528 13125 19552
rect 12805 18464 12813 18528
rect 12877 18464 12893 18528
rect 12957 18464 12973 18528
rect 13037 18464 13053 18528
rect 13117 18464 13125 18528
rect 12805 17440 13125 18464
rect 12805 17376 12813 17440
rect 12877 17376 12893 17440
rect 12957 17376 12973 17440
rect 13037 17376 13053 17440
rect 13117 17376 13125 17440
rect 12805 16352 13125 17376
rect 12805 16288 12813 16352
rect 12877 16288 12893 16352
rect 12957 16288 12973 16352
rect 13037 16288 13053 16352
rect 13117 16288 13125 16352
rect 12805 15264 13125 16288
rect 12805 15200 12813 15264
rect 12877 15200 12893 15264
rect 12957 15200 12973 15264
rect 13037 15200 13053 15264
rect 13117 15200 13125 15264
rect 12805 14176 13125 15200
rect 12805 14112 12813 14176
rect 12877 14112 12893 14176
rect 12957 14112 12973 14176
rect 13037 14112 13053 14176
rect 13117 14112 13125 14176
rect 12805 13088 13125 14112
rect 12805 13024 12813 13088
rect 12877 13024 12893 13088
rect 12957 13024 12973 13088
rect 13037 13024 13053 13088
rect 13117 13024 13125 13088
rect 12805 12000 13125 13024
rect 12805 11936 12813 12000
rect 12877 11936 12893 12000
rect 12957 11936 12973 12000
rect 13037 11936 13053 12000
rect 13117 11936 13125 12000
rect 12805 10912 13125 11936
rect 12805 10848 12813 10912
rect 12877 10848 12893 10912
rect 12957 10848 12973 10912
rect 13037 10848 13053 10912
rect 13117 10848 13125 10912
rect 12805 9824 13125 10848
rect 12805 9760 12813 9824
rect 12877 9760 12893 9824
rect 12957 9760 12973 9824
rect 13037 9760 13053 9824
rect 13117 9760 13125 9824
rect 12805 8736 13125 9760
rect 12805 8672 12813 8736
rect 12877 8672 12893 8736
rect 12957 8672 12973 8736
rect 13037 8672 13053 8736
rect 13117 8672 13125 8736
rect 12805 7648 13125 8672
rect 12805 7584 12813 7648
rect 12877 7584 12893 7648
rect 12957 7584 12973 7648
rect 13037 7584 13053 7648
rect 13117 7584 13125 7648
rect 12805 6560 13125 7584
rect 12805 6496 12813 6560
rect 12877 6496 12893 6560
rect 12957 6496 12973 6560
rect 13037 6496 13053 6560
rect 13117 6496 13125 6560
rect 12805 5472 13125 6496
rect 12805 5408 12813 5472
rect 12877 5408 12893 5472
rect 12957 5408 12973 5472
rect 13037 5408 13053 5472
rect 13117 5408 13125 5472
rect 12805 4384 13125 5408
rect 12805 4320 12813 4384
rect 12877 4320 12893 4384
rect 12957 4320 12973 4384
rect 13037 4320 13053 4384
rect 13117 4320 13125 4384
rect 12805 3296 13125 4320
rect 12805 3232 12813 3296
rect 12877 3232 12893 3296
rect 12957 3232 12973 3296
rect 13037 3232 13053 3296
rect 13117 3232 13125 3296
rect 12805 2208 13125 3232
rect 12805 2144 12813 2208
rect 12877 2144 12893 2208
rect 12957 2144 12973 2208
rect 13037 2144 13053 2208
rect 13117 2144 13125 2208
rect 12805 2128 13125 2144
rect 15770 24512 16091 25536
rect 15770 24448 15778 24512
rect 15842 24448 15858 24512
rect 15922 24448 15938 24512
rect 16002 24448 16018 24512
rect 16082 24448 16091 24512
rect 15770 23424 16091 24448
rect 15770 23360 15778 23424
rect 15842 23360 15858 23424
rect 15922 23360 15938 23424
rect 16002 23360 16018 23424
rect 16082 23360 16091 23424
rect 15770 22336 16091 23360
rect 15770 22272 15778 22336
rect 15842 22272 15858 22336
rect 15922 22272 15938 22336
rect 16002 22272 16018 22336
rect 16082 22272 16091 22336
rect 15770 21248 16091 22272
rect 15770 21184 15778 21248
rect 15842 21184 15858 21248
rect 15922 21184 15938 21248
rect 16002 21184 16018 21248
rect 16082 21184 16091 21248
rect 15770 20160 16091 21184
rect 15770 20096 15778 20160
rect 15842 20096 15858 20160
rect 15922 20096 15938 20160
rect 16002 20096 16018 20160
rect 16082 20096 16091 20160
rect 15770 19072 16091 20096
rect 15770 19008 15778 19072
rect 15842 19008 15858 19072
rect 15922 19008 15938 19072
rect 16002 19008 16018 19072
rect 16082 19008 16091 19072
rect 15770 17984 16091 19008
rect 15770 17920 15778 17984
rect 15842 17920 15858 17984
rect 15922 17920 15938 17984
rect 16002 17920 16018 17984
rect 16082 17920 16091 17984
rect 15770 16896 16091 17920
rect 15770 16832 15778 16896
rect 15842 16832 15858 16896
rect 15922 16832 15938 16896
rect 16002 16832 16018 16896
rect 16082 16832 16091 16896
rect 15770 15808 16091 16832
rect 15770 15744 15778 15808
rect 15842 15744 15858 15808
rect 15922 15744 15938 15808
rect 16002 15744 16018 15808
rect 16082 15744 16091 15808
rect 15770 14720 16091 15744
rect 15770 14656 15778 14720
rect 15842 14656 15858 14720
rect 15922 14656 15938 14720
rect 16002 14656 16018 14720
rect 16082 14656 16091 14720
rect 15770 13632 16091 14656
rect 15770 13568 15778 13632
rect 15842 13568 15858 13632
rect 15922 13568 15938 13632
rect 16002 13568 16018 13632
rect 16082 13568 16091 13632
rect 15770 12544 16091 13568
rect 15770 12480 15778 12544
rect 15842 12480 15858 12544
rect 15922 12480 15938 12544
rect 16002 12480 16018 12544
rect 16082 12480 16091 12544
rect 15770 11456 16091 12480
rect 15770 11392 15778 11456
rect 15842 11392 15858 11456
rect 15922 11392 15938 11456
rect 16002 11392 16018 11456
rect 16082 11392 16091 11456
rect 15770 10368 16091 11392
rect 15770 10304 15778 10368
rect 15842 10304 15858 10368
rect 15922 10304 15938 10368
rect 16002 10304 16018 10368
rect 16082 10304 16091 10368
rect 15770 9280 16091 10304
rect 15770 9216 15778 9280
rect 15842 9216 15858 9280
rect 15922 9216 15938 9280
rect 16002 9216 16018 9280
rect 16082 9216 16091 9280
rect 15770 8192 16091 9216
rect 15770 8128 15778 8192
rect 15842 8128 15858 8192
rect 15922 8128 15938 8192
rect 16002 8128 16018 8192
rect 16082 8128 16091 8192
rect 15770 7104 16091 8128
rect 15770 7040 15778 7104
rect 15842 7040 15858 7104
rect 15922 7040 15938 7104
rect 16002 7040 16018 7104
rect 16082 7040 16091 7104
rect 15770 6016 16091 7040
rect 15770 5952 15778 6016
rect 15842 5952 15858 6016
rect 15922 5952 15938 6016
rect 16002 5952 16018 6016
rect 16082 5952 16091 6016
rect 15770 4928 16091 5952
rect 15770 4864 15778 4928
rect 15842 4864 15858 4928
rect 15922 4864 15938 4928
rect 16002 4864 16018 4928
rect 16082 4864 16091 4928
rect 15770 3840 16091 4864
rect 15770 3776 15778 3840
rect 15842 3776 15858 3840
rect 15922 3776 15938 3840
rect 16002 3776 16018 3840
rect 16082 3776 16091 3840
rect 15770 2752 16091 3776
rect 16622 2957 16682 33219
rect 16619 2956 16685 2957
rect 16619 2892 16620 2956
rect 16684 2892 16685 2956
rect 16619 2891 16685 2892
rect 15770 2688 15778 2752
rect 15842 2688 15858 2752
rect 15922 2688 15938 2752
rect 16002 2688 16018 2752
rect 16082 2688 16091 2752
rect 15770 2128 16091 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__051__B asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__B
timestamp 1644511149
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__A1
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__A
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__A
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1644511149
transform 1 0 13432 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B
timestamp 1644511149
transform -1 0 13708 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__B
timestamp 1644511149
transform 1 0 16008 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__B
timestamp 1644511149
transform 1 0 12880 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A2
timestamp 1644511149
transform -1 0 13708 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__C1
timestamp 1644511149
transform -1 0 12788 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A2
timestamp 1644511149
transform -1 0 17204 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1644511149
transform -1 0 14628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 1564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 1564 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 18124 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 1748 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 17112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 16192 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 15732 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 1564 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 15548 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 16836 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 16928 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 2208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 17572 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 17480 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 17480 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 17572 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 17572 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 13616 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1644511149
transform -1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output25_A
timestamp 1644511149
transform -1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output29_A
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1644511149
transform 1 0 2024 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22
timestamp 1644511149
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1644511149
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1644511149
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_128
timestamp 1644511149
transform 1 0 12880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1644511149
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_182 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_13
timestamp 1644511149
transform 1 0 2300 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_25
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_37
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1644511149
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_181
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_186
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1644511149
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp 1644511149
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1644511149
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_189
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_7
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_23
timestamp 1644511149
transform 1 0 3220 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_35
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1644511149
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1644511149
transform 1 0 17204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1644511149
transform 1 0 17480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1644511149
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1644511149
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1644511149
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_5
timestamp 1644511149
transform 1 0 1564 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_17
timestamp 1644511149
transform 1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1644511149
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_13
timestamp 1644511149
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_25
timestamp 1644511149
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_37
timestamp 1644511149
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1644511149
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_183
timestamp 1644511149
transform 1 0 17940 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_186
timestamp 1644511149
transform 1 0 18216 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1644511149
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_186
timestamp 1644511149
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_113
timestamp 1644511149
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_125
timestamp 1644511149
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1644511149
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_101
timestamp 1644511149
transform 1 0 10396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_118
timestamp 1644511149
transform 1 0 11960 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_130
timestamp 1644511149
transform 1 0 13064 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_142
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1644511149
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1644511149
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_5
timestamp 1644511149
transform 1 0 1564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1644511149
transform 1 0 2668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1644511149
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1644511149
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1644511149
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_147
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_189
timestamp 1644511149
transform 1 0 18492 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_13
timestamp 1644511149
transform 1 0 2300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1644511149
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_131
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1644511149
transform 1 0 14628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_159
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_189
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_127
timestamp 1644511149
transform 1 0 12788 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_143
timestamp 1644511149
transform 1 0 14260 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_155
timestamp 1644511149
transform 1 0 15364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_167
timestamp 1644511149
transform 1 0 16468 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_175
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1644511149
transform 1 0 17572 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_186
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_189
timestamp 1644511149
transform 1 0 18492 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_116
timestamp 1644511149
transform 1 0 11776 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_130
timestamp 1644511149
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_189
timestamp 1644511149
transform 1 0 18492 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_7
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1644511149
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_129
timestamp 1644511149
transform 1 0 12972 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_132
timestamp 1644511149
transform 1 0 13248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_145
timestamp 1644511149
transform 1 0 14444 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_157
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1644511149
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_189
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_189
timestamp 1644511149
transform 1 0 18492 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_189
timestamp 1644511149
transform 1 0 18492 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_179
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_186
timestamp 1644511149
transform 1 0 18216 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_189
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_159
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_163
timestamp 1644511149
transform 1 0 16100 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_175
timestamp 1644511149
transform 1 0 17204 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1644511149
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_5
timestamp 1644511149
transform 1 0 1564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_17
timestamp 1644511149
transform 1 0 2668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_29
timestamp 1644511149
transform 1 0 3772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_41
timestamp 1644511149
transform 1 0 4876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1644511149
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_157
timestamp 1644511149
transform 1 0 15548 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_172
timestamp 1644511149
transform 1 0 16928 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_179
timestamp 1644511149
transform 1 0 17572 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_186
timestamp 1644511149
transform 1 0 18216 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_13
timestamp 1644511149
transform 1 0 2300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_25
timestamp 1644511149
transform 1 0 3404 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_159
timestamp 1644511149
transform 1 0 15732 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_163
timestamp 1644511149
transform 1 0 16100 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_172
timestamp 1644511149
transform 1 0 16928 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_181
timestamp 1644511149
transform 1 0 17756 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_158
timestamp 1644511149
transform 1 0 15640 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_175
timestamp 1644511149
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_184
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_143
timestamp 1644511149
transform 1 0 14260 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_147
timestamp 1644511149
transform 1 0 14628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_170
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_181
timestamp 1644511149
transform 1 0 17756 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_133
timestamp 1644511149
transform 1 0 13340 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_144
timestamp 1644511149
transform 1 0 14352 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_154
timestamp 1644511149
transform 1 0 15272 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_178
timestamp 1644511149
transform 1 0 17480 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_185
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_189
timestamp 1644511149
transform 1 0 18492 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_127
timestamp 1644511149
transform 1 0 12788 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_130
timestamp 1644511149
transform 1 0 13064 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_147
timestamp 1644511149
transform 1 0 14628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_151
timestamp 1644511149
transform 1 0 14996 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_159
timestamp 1644511149
transform 1 0 15732 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_184
timestamp 1644511149
transform 1 0 18032 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_130
timestamp 1644511149
transform 1 0 13064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_139
timestamp 1644511149
transform 1 0 13892 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_148
timestamp 1644511149
transform 1 0 14720 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_186
timestamp 1644511149
transform 1 0 18216 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_127
timestamp 1644511149
transform 1 0 12788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_150
timestamp 1644511149
transform 1 0 14904 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_161
timestamp 1644511149
transform 1 0 15916 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_178
timestamp 1644511149
transform 1 0 17480 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_186
timestamp 1644511149
transform 1 0 18216 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_133
timestamp 1644511149
transform 1 0 13340 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_144
timestamp 1644511149
transform 1 0 14352 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_153
timestamp 1644511149
transform 1 0 15180 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_173
timestamp 1644511149
transform 1 0 17020 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_185
timestamp 1644511149
transform 1 0 18124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_189
timestamp 1644511149
transform 1 0 18492 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_157
timestamp 1644511149
transform 1 0 15548 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_183
timestamp 1644511149
transform 1 0 17940 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_7
timestamp 1644511149
transform 1 0 1748 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_19
timestamp 1644511149
transform 1 0 2852 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_31
timestamp 1644511149
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_43
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_153
timestamp 1644511149
transform 1 0 15180 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_157
timestamp 1644511149
transform 1 0 15548 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_172
timestamp 1644511149
transform 1 0 16928 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_183
timestamp 1644511149
transform 1 0 17940 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_189
timestamp 1644511149
transform 1 0 18492 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_11
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1644511149
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_159
timestamp 1644511149
transform 1 0 15732 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_170
timestamp 1644511149
transform 1 0 16744 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_178
timestamp 1644511149
transform 1 0 17480 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_186
timestamp 1644511149
transform 1 0 18216 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_173
timestamp 1644511149
transform 1 0 17020 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_177
timestamp 1644511149
transform 1 0 17388 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_186
timestamp 1644511149
transform 1 0 18216 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1644511149
transform 1 0 17204 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_186
timestamp 1644511149
transform 1 0 18216 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_189
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_189
timestamp 1644511149
transform 1 0 18492 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_189
timestamp 1644511149
transform 1 0 18492 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_179
timestamp 1644511149
transform 1 0 17572 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_186
timestamp 1644511149
transform 1 0 18216 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_13
timestamp 1644511149
transform 1 0 2300 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_25
timestamp 1644511149
transform 1 0 3404 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_37
timestamp 1644511149
transform 1 0 4508 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1644511149
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_189
timestamp 1644511149
transform 1 0 18492 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_189
timestamp 1644511149
transform 1 0 18492 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_175
timestamp 1644511149
transform 1 0 17204 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_178
timestamp 1644511149
transform 1 0 17480 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_186
timestamp 1644511149
transform 1 0 18216 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_169
timestamp 1644511149
transform 1 0 16652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_172
timestamp 1644511149
transform 1 0 16928 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_178
timestamp 1644511149
transform 1 0 17480 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_186
timestamp 1644511149
transform 1 0 18216 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1644511149
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_173
timestamp 1644511149
transform 1 0 17020 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_178
timestamp 1644511149
transform 1 0 17480 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_186
timestamp 1644511149
transform 1 0 18216 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_6
timestamp 1644511149
transform 1 0 1656 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_12
timestamp 1644511149
transform 1 0 2208 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_144
timestamp 1644511149
transform 1 0 14352 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_151
timestamp 1644511149
transform 1 0 14996 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_157
timestamp 1644511149
transform 1 0 15548 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_163
timestamp 1644511149
transform 1 0 16100 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_168
timestamp 1644511149
transform 1 0 16560 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_182
timestamp 1644511149
transform 1 0 17848 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_6
timestamp 1644511149
transform 1 0 1656 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_13
timestamp 1644511149
transform 1 0 2300 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_20
timestamp 1644511149
transform 1 0 2944 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_29
timestamp 1644511149
transform 1 0 3772 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_44
timestamp 1644511149
transform 1 0 5152 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_64
timestamp 1644511149
transform 1 0 6992 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_70
timestamp 1644511149
transform 1 0 7544 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_74
timestamp 1644511149
transform 1 0 7912 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_80
timestamp 1644511149
transform 1 0 8464 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_84
timestamp 1644511149
transform 1 0 8832 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_90
timestamp 1644511149
transform 1 0 9384 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_94
timestamp 1644511149
transform 1 0 9752 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_120
timestamp 1644511149
transform 1 0 12144 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_126
timestamp 1644511149
transform 1 0 12696 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_130
timestamp 1644511149
transform 1 0 13064 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_141
timestamp 1644511149
transform 1 0 14076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_145
timestamp 1644511149
transform 1 0 14444 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_153
timestamp 1644511149
transform 1 0 15180 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_171
timestamp 1644511149
transform 1 0 16836 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_175
timestamp 1644511149
transform 1 0 17204 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_186
timestamp 1644511149
transform 1 0 18216 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_7
timestamp 1644511149
transform 1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_14
timestamp 1644511149
transform 1 0 2392 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1644511149
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_32
timestamp 1644511149
transform 1 0 4048 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_39
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_46
timestamp 1644511149
transform 1 0 5336 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_54
timestamp 1644511149
transform 1 0 6072 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_60
timestamp 1644511149
transform 1 0 6624 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_67
timestamp 1644511149
transform 1 0 7268 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_74
timestamp 1644511149
transform 1 0 7912 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_82
timestamp 1644511149
transform 1 0 8648 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_88
timestamp 1644511149
transform 1 0 9200 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_95
timestamp 1644511149
transform 1 0 9844 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_102
timestamp 1644511149
transform 1 0 10488 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_110
timestamp 1644511149
transform 1 0 11224 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_116
timestamp 1644511149
transform 1 0 11776 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_123
timestamp 1644511149
transform 1 0 12420 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_130
timestamp 1644511149
transform 1 0 13064 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1644511149
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_145
timestamp 1644511149
transform 1 0 14444 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_150
timestamp 1644511149
transform 1 0 14904 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_164
timestamp 1644511149
transform 1 0 16192 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_179
timestamp 1644511149
transform 1 0 17572 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_185
timestamp 1644511149
transform 1 0 18124 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 18860 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 18860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 18860 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 18860 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 18860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 18860 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 18860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _046_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18216 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _047_
timestamp 1644511149
transform -1 0 14904 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _048_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _049_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _050_
timestamp 1644511149
transform 1 0 15824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _051_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _052_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _053_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _054_
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _055_
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _056_
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _057_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _058_
timestamp 1644511149
transform -1 0 16928 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _059_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _060_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _061_
timestamp 1644511149
transform 1 0 14260 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _062_
timestamp 1644511149
transform -1 0 16744 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_4  _063_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16100 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _064_
timestamp 1644511149
transform 1 0 17940 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _065_
timestamp 1644511149
transform -1 0 17572 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _066_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _067_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _068_
timestamp 1644511149
transform 1 0 17848 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _069_
timestamp 1644511149
transform 1 0 13432 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _070_
timestamp 1644511149
transform 1 0 14720 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _071_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _072_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17480 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _073_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16192 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _074_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _075_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 18216 0 -1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _076_
timestamp 1644511149
transform -1 0 16192 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _077_
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _078_
timestamp 1644511149
transform -1 0 18216 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _079_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _080_
timestamp 1644511149
transform -1 0 13524 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _081_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _082_
timestamp 1644511149
transform -1 0 13708 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _083_
timestamp 1644511149
transform -1 0 11776 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _084_
timestamp 1644511149
transform -1 0 16100 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _085_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _086_
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _087_
timestamp 1644511149
transform -1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _088_
timestamp 1644511149
transform 1 0 15548 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _089_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _090_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 15272 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1644511149
transform 1 0 16468 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _092_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _093_
timestamp 1644511149
transform 1 0 17296 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _094_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16744 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__a31o_1  _095_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _096_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 15548 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _097_ asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _098_
timestamp 1644511149
transform -1 0 17940 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _099_
timestamp 1644511149
transform -1 0 13616 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _100_
timestamp 1644511149
transform -1 0 17940 0 1 34816
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _101_
timestamp 1644511149
transform 1 0 14076 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _102_
timestamp 1644511149
transform 1 0 17572 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  _103__44 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _104__45
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _105__46
timestamp 1644511149
transform 1 0 2116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _106__47
timestamp 1644511149
transform 1 0 2024 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _107__48
timestamp 1644511149
transform 1 0 2760 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _108__49
timestamp 1644511149
transform 1 0 2668 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _109__50
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _110__51
timestamp 1644511149
transform 1 0 3496 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _111__52
timestamp 1644511149
transform 1 0 4416 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _112__53
timestamp 1644511149
transform 1 0 5060 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _113__54
timestamp 1644511149
transform 1 0 4876 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _114__55
timestamp 1644511149
transform 1 0 5520 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _115__56
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _116__57
timestamp 1644511149
transform 1 0 6992 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _117__58
timestamp 1644511149
transform 1 0 6716 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _118__59
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _119__60
timestamp 1644511149
transform 1 0 7636 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _120__61
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _121__62
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _122__63
timestamp 1644511149
transform 1 0 9568 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _123__64
timestamp 1644511149
transform 1 0 14168 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _124__33
timestamp 1644511149
transform -1 0 9752 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _125__34
timestamp 1644511149
transform -1 0 10488 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _126__35
timestamp 1644511149
transform -1 0 10764 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _127__36
timestamp 1644511149
transform -1 0 11776 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _128__37
timestamp 1644511149
transform -1 0 12420 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _129__38
timestamp 1644511149
transform -1 0 12144 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _130__39
timestamp 1644511149
transform -1 0 13064 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _131__40
timestamp 1644511149
transform -1 0 13064 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _132__41
timestamp 1644511149
transform -1 0 13708 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _133__42
timestamp 1644511149
transform -1 0 14352 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _134__43
timestamp 1644511149
transform -1 0 14996 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform -1 0 18216 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input7 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1644511149
transform 1 0 17296 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform -1 0 15548 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1644511149
transform -1 0 15916 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1644511149
transform -1 0 16192 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1644511149
transform 1 0 16928 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input15 asic/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 17940 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform -1 0 18216 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1644511149
transform -1 0 18216 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 17940 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1644511149
transform -1 0 14904 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1644511149
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1644511149
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1644511149
transform -1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1644511149
transform 1 0 17112 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1644511149
transform -1 0 16560 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1644511149
transform -1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1644511149
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1644511149
transform -1 0 15180 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1644511149
transform -1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1644511149
transform -1 0 18216 0 -1 44608
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 8168 800 8288 6 A[0]
port 0 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 A[1]
port 1 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 A[2]
port 2 nsew signal input
rlabel metal2 s 16394 49200 16450 50000 6 A[3]
port 3 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 A[4]
port 4 nsew signal input
rlabel metal3 s 19200 15648 20000 15768 6 A[5]
port 5 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 A[6]
port 6 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 A[7]
port 7 nsew signal input
rlabel metal2 s 19614 49200 19670 50000 6 A[8]
port 8 nsew signal input
rlabel metal3 s 19200 34416 20000 34536 6 A[9]
port 9 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 B[0]
port 10 nsew signal input
rlabel metal2 s 15474 49200 15530 50000 6 B[1]
port 11 nsew signal input
rlabel metal2 s 15934 49200 15990 50000 6 B[2]
port 12 nsew signal input
rlabel metal2 s 16854 49200 16910 50000 6 B[3]
port 13 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 B[4]
port 14 nsew signal input
rlabel metal3 s 19200 21904 20000 22024 6 B[5]
port 15 nsew signal input
rlabel metal2 s 18234 49200 18290 50000 6 B[6]
port 16 nsew signal input
rlabel metal2 s 18694 49200 18750 50000 6 B[7]
port 17 nsew signal input
rlabel metal3 s 19200 28160 20000 28280 6 B[8]
port 18 nsew signal input
rlabel metal3 s 19200 40672 20000 40792 6 B[9]
port 19 nsew signal input
rlabel metal2 s 15014 49200 15070 50000 6 Ci
port 20 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 Co
port 21 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 S[0]
port 22 nsew signal tristate
rlabel metal3 s 0 24896 800 25016 6 S[1]
port 23 nsew signal tristate
rlabel metal3 s 19200 9392 20000 9512 6 S[2]
port 24 nsew signal tristate
rlabel metal2 s 17314 49200 17370 50000 6 S[3]
port 25 nsew signal tristate
rlabel metal2 s 17774 49200 17830 50000 6 S[4]
port 26 nsew signal tristate
rlabel metal2 s 7470 0 7526 800 6 S[5]
port 27 nsew signal tristate
rlabel metal3 s 0 41624 800 41744 6 S[6]
port 28 nsew signal tristate
rlabel metal2 s 19154 49200 19210 50000 6 S[7]
port 29 nsew signal tristate
rlabel metal3 s 0 47200 800 47320 6 S[8]
port 30 nsew signal tristate
rlabel metal3 s 19200 46928 20000 47048 6 S[9]
port 31 nsew signal tristate
rlabel metal2 s 202 49200 258 50000 6 io_oeb[0]
port 32 nsew signal tristate
rlabel metal2 s 4802 49200 4858 50000 6 io_oeb[10]
port 33 nsew signal tristate
rlabel metal2 s 5262 49200 5318 50000 6 io_oeb[11]
port 34 nsew signal tristate
rlabel metal2 s 5722 49200 5778 50000 6 io_oeb[12]
port 35 nsew signal tristate
rlabel metal2 s 6182 49200 6238 50000 6 io_oeb[13]
port 36 nsew signal tristate
rlabel metal2 s 6642 49200 6698 50000 6 io_oeb[14]
port 37 nsew signal tristate
rlabel metal2 s 7102 49200 7158 50000 6 io_oeb[15]
port 38 nsew signal tristate
rlabel metal2 s 7562 49200 7618 50000 6 io_oeb[16]
port 39 nsew signal tristate
rlabel metal2 s 8022 49200 8078 50000 6 io_oeb[17]
port 40 nsew signal tristate
rlabel metal2 s 8482 49200 8538 50000 6 io_oeb[18]
port 41 nsew signal tristate
rlabel metal2 s 8942 49200 8998 50000 6 io_oeb[19]
port 42 nsew signal tristate
rlabel metal2 s 662 49200 718 50000 6 io_oeb[1]
port 43 nsew signal tristate
rlabel metal2 s 9402 49200 9458 50000 6 io_oeb[20]
port 44 nsew signal tristate
rlabel metal2 s 9862 49200 9918 50000 6 io_oeb[21]
port 45 nsew signal tristate
rlabel metal2 s 10414 49200 10470 50000 6 io_oeb[22]
port 46 nsew signal tristate
rlabel metal2 s 10874 49200 10930 50000 6 io_oeb[23]
port 47 nsew signal tristate
rlabel metal2 s 11334 49200 11390 50000 6 io_oeb[24]
port 48 nsew signal tristate
rlabel metal2 s 11794 49200 11850 50000 6 io_oeb[25]
port 49 nsew signal tristate
rlabel metal2 s 12254 49200 12310 50000 6 io_oeb[26]
port 50 nsew signal tristate
rlabel metal2 s 12714 49200 12770 50000 6 io_oeb[27]
port 51 nsew signal tristate
rlabel metal2 s 13174 49200 13230 50000 6 io_oeb[28]
port 52 nsew signal tristate
rlabel metal2 s 13634 49200 13690 50000 6 io_oeb[29]
port 53 nsew signal tristate
rlabel metal2 s 1122 49200 1178 50000 6 io_oeb[2]
port 54 nsew signal tristate
rlabel metal2 s 14094 49200 14150 50000 6 io_oeb[30]
port 55 nsew signal tristate
rlabel metal2 s 14554 49200 14610 50000 6 io_oeb[31]
port 56 nsew signal tristate
rlabel metal2 s 1582 49200 1638 50000 6 io_oeb[3]
port 57 nsew signal tristate
rlabel metal2 s 2042 49200 2098 50000 6 io_oeb[4]
port 58 nsew signal tristate
rlabel metal2 s 2502 49200 2558 50000 6 io_oeb[5]
port 59 nsew signal tristate
rlabel metal2 s 2962 49200 3018 50000 6 io_oeb[6]
port 60 nsew signal tristate
rlabel metal2 s 3422 49200 3478 50000 6 io_oeb[7]
port 61 nsew signal tristate
rlabel metal2 s 3882 49200 3938 50000 6 io_oeb[8]
port 62 nsew signal tristate
rlabel metal2 s 4342 49200 4398 50000 6 io_oeb[9]
port 63 nsew signal tristate
rlabel metal4 s 3910 2128 4230 47376 6 vccd1
port 64 nsew power input
rlabel metal4 s 9840 2128 10160 47376 6 vccd1
port 64 nsew power input
rlabel metal4 s 15771 2128 16091 47376 6 vccd1
port 64 nsew power input
rlabel metal4 s 6874 2128 7194 47376 6 vssd1
port 65 nsew ground input
rlabel metal4 s 12805 2128 13125 47376 6 vssd1
port 65 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 20000 50000
<< end >>

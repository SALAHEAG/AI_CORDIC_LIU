magic
tech sky130A
magscale 1 2
timestamp 1695401851
<< obsli1 >>
rect 1104 2159 18860 47345
<< obsm1 >>
rect 198 2128 19674 47456
<< metal2 >>
rect 202 49200 258 50000
rect 662 49200 718 50000
rect 1122 49200 1178 50000
rect 1582 49200 1638 50000
rect 2042 49200 2098 50000
rect 2502 49200 2558 50000
rect 2962 49200 3018 50000
rect 3422 49200 3478 50000
rect 3882 49200 3938 50000
rect 4342 49200 4398 50000
rect 4802 49200 4858 50000
rect 5262 49200 5318 50000
rect 5722 49200 5778 50000
rect 6182 49200 6238 50000
rect 6642 49200 6698 50000
rect 7102 49200 7158 50000
rect 7562 49200 7618 50000
rect 8022 49200 8078 50000
rect 8482 49200 8538 50000
rect 8942 49200 8998 50000
rect 9402 49200 9458 50000
rect 9862 49200 9918 50000
rect 10414 49200 10470 50000
rect 10874 49200 10930 50000
rect 11334 49200 11390 50000
rect 11794 49200 11850 50000
rect 12254 49200 12310 50000
rect 12714 49200 12770 50000
rect 13174 49200 13230 50000
rect 13634 49200 13690 50000
rect 14094 49200 14150 50000
rect 14554 49200 14610 50000
rect 15014 49200 15070 50000
rect 15474 49200 15530 50000
rect 15934 49200 15990 50000
rect 16394 49200 16450 50000
rect 16854 49200 16910 50000
rect 17314 49200 17370 50000
rect 17774 49200 17830 50000
rect 18234 49200 18290 50000
rect 18694 49200 18750 50000
rect 19154 49200 19210 50000
rect 19614 49200 19670 50000
rect 2502 0 2558 800
rect 7470 0 7526 800
rect 12438 0 12494 800
rect 17406 0 17462 800
<< obsm2 >>
rect 314 49144 606 49314
rect 774 49144 1066 49314
rect 1234 49144 1526 49314
rect 1694 49144 1986 49314
rect 2154 49144 2446 49314
rect 2614 49144 2906 49314
rect 3074 49144 3366 49314
rect 3534 49144 3826 49314
rect 3994 49144 4286 49314
rect 4454 49144 4746 49314
rect 4914 49144 5206 49314
rect 5374 49144 5666 49314
rect 5834 49144 6126 49314
rect 6294 49144 6586 49314
rect 6754 49144 7046 49314
rect 7214 49144 7506 49314
rect 7674 49144 7966 49314
rect 8134 49144 8426 49314
rect 8594 49144 8886 49314
rect 9054 49144 9346 49314
rect 9514 49144 9806 49314
rect 9974 49144 10358 49314
rect 10526 49144 10818 49314
rect 10986 49144 11278 49314
rect 11446 49144 11738 49314
rect 11906 49144 12198 49314
rect 12366 49144 12658 49314
rect 12826 49144 13118 49314
rect 13286 49144 13578 49314
rect 13746 49144 14038 49314
rect 14206 49144 14498 49314
rect 14666 49144 14958 49314
rect 15126 49144 15418 49314
rect 15586 49144 15878 49314
rect 16046 49144 16338 49314
rect 16506 49144 16798 49314
rect 16966 49144 17258 49314
rect 17426 49144 17718 49314
rect 17886 49144 18178 49314
rect 18346 49144 18638 49314
rect 18806 49144 19098 49314
rect 19266 49144 19558 49314
rect 204 856 19668 49144
rect 204 800 2446 856
rect 2614 800 7414 856
rect 7582 800 12382 856
rect 12550 800 17350 856
rect 17518 800 19668 856
<< metal3 >>
rect 0 47200 800 47320
rect 19200 46928 20000 47048
rect 0 41624 800 41744
rect 19200 40672 20000 40792
rect 0 36048 800 36168
rect 19200 34416 20000 34536
rect 0 30472 800 30592
rect 19200 28160 20000 28280
rect 0 24896 800 25016
rect 19200 21904 20000 22024
rect 0 19320 800 19440
rect 19200 15648 20000 15768
rect 0 13744 800 13864
rect 19200 9392 20000 9512
rect 0 8168 800 8288
rect 19200 3136 20000 3256
rect 0 2728 800 2848
<< obsm3 >>
rect 880 47128 19200 47361
rect 880 47120 19120 47128
rect 800 46848 19120 47120
rect 800 41824 19200 46848
rect 880 41544 19200 41824
rect 800 40872 19200 41544
rect 800 40592 19120 40872
rect 800 36248 19200 40592
rect 880 35968 19200 36248
rect 800 34616 19200 35968
rect 800 34336 19120 34616
rect 800 30672 19200 34336
rect 880 30392 19200 30672
rect 800 28360 19200 30392
rect 800 28080 19120 28360
rect 800 25096 19200 28080
rect 880 24816 19200 25096
rect 800 22104 19200 24816
rect 800 21824 19120 22104
rect 800 19520 19200 21824
rect 880 19240 19200 19520
rect 800 15848 19200 19240
rect 800 15568 19120 15848
rect 800 13944 19200 15568
rect 880 13664 19200 13944
rect 800 9592 19200 13664
rect 800 9312 19120 9592
rect 800 8368 19200 9312
rect 880 8088 19200 8368
rect 800 3336 19200 8088
rect 800 3056 19120 3336
rect 800 2928 19200 3056
rect 880 2648 19200 2928
rect 800 2143 19200 2648
<< metal4 >>
rect 3910 2128 4230 47376
rect 6874 2128 7194 47376
rect 9840 2128 10160 47376
rect 12805 2128 13125 47376
rect 15771 2128 16091 47376
<< obsm4 >>
rect 4310 2128 6794 47376
rect 7274 2128 9760 47376
rect 10240 2128 12725 47376
rect 13205 2128 15691 47376
rect 16171 2128 16685 47376
<< labels >>
rlabel metal3 s 0 8168 800 8288 6 A[0]
port 1 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 A[2]
port 3 nsew signal input
rlabel metal2 s 16394 49200 16450 50000 6 A[3]
port 4 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 A[4]
port 5 nsew signal input
rlabel metal3 s 19200 15648 20000 15768 6 A[5]
port 6 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 A[6]
port 7 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 A[7]
port 8 nsew signal input
rlabel metal2 s 19614 49200 19670 50000 6 A[8]
port 9 nsew signal input
rlabel metal3 s 19200 34416 20000 34536 6 A[9]
port 10 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 B[0]
port 11 nsew signal input
rlabel metal2 s 15474 49200 15530 50000 6 B[1]
port 12 nsew signal input
rlabel metal2 s 15934 49200 15990 50000 6 B[2]
port 13 nsew signal input
rlabel metal2 s 16854 49200 16910 50000 6 B[3]
port 14 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 B[4]
port 15 nsew signal input
rlabel metal3 s 19200 21904 20000 22024 6 B[5]
port 16 nsew signal input
rlabel metal2 s 18234 49200 18290 50000 6 B[6]
port 17 nsew signal input
rlabel metal2 s 18694 49200 18750 50000 6 B[7]
port 18 nsew signal input
rlabel metal3 s 19200 28160 20000 28280 6 B[8]
port 19 nsew signal input
rlabel metal3 s 19200 40672 20000 40792 6 B[9]
port 20 nsew signal input
rlabel metal2 s 15014 49200 15070 50000 6 Ci
port 21 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 Co
port 22 nsew signal output
rlabel metal3 s 19200 3136 20000 3256 6 S[0]
port 23 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 S[1]
port 24 nsew signal output
rlabel metal3 s 19200 9392 20000 9512 6 S[2]
port 25 nsew signal output
rlabel metal2 s 17314 49200 17370 50000 6 S[3]
port 26 nsew signal output
rlabel metal2 s 17774 49200 17830 50000 6 S[4]
port 27 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 S[5]
port 28 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 S[6]
port 29 nsew signal output
rlabel metal2 s 19154 49200 19210 50000 6 S[7]
port 30 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 S[8]
port 31 nsew signal output
rlabel metal3 s 19200 46928 20000 47048 6 S[9]
port 32 nsew signal output
rlabel metal2 s 202 49200 258 50000 6 io_oeb[0]
port 33 nsew signal output
rlabel metal2 s 4802 49200 4858 50000 6 io_oeb[10]
port 34 nsew signal output
rlabel metal2 s 5262 49200 5318 50000 6 io_oeb[11]
port 35 nsew signal output
rlabel metal2 s 5722 49200 5778 50000 6 io_oeb[12]
port 36 nsew signal output
rlabel metal2 s 6182 49200 6238 50000 6 io_oeb[13]
port 37 nsew signal output
rlabel metal2 s 6642 49200 6698 50000 6 io_oeb[14]
port 38 nsew signal output
rlabel metal2 s 7102 49200 7158 50000 6 io_oeb[15]
port 39 nsew signal output
rlabel metal2 s 7562 49200 7618 50000 6 io_oeb[16]
port 40 nsew signal output
rlabel metal2 s 8022 49200 8078 50000 6 io_oeb[17]
port 41 nsew signal output
rlabel metal2 s 8482 49200 8538 50000 6 io_oeb[18]
port 42 nsew signal output
rlabel metal2 s 8942 49200 8998 50000 6 io_oeb[19]
port 43 nsew signal output
rlabel metal2 s 662 49200 718 50000 6 io_oeb[1]
port 44 nsew signal output
rlabel metal2 s 9402 49200 9458 50000 6 io_oeb[20]
port 45 nsew signal output
rlabel metal2 s 9862 49200 9918 50000 6 io_oeb[21]
port 46 nsew signal output
rlabel metal2 s 10414 49200 10470 50000 6 io_oeb[22]
port 47 nsew signal output
rlabel metal2 s 10874 49200 10930 50000 6 io_oeb[23]
port 48 nsew signal output
rlabel metal2 s 11334 49200 11390 50000 6 io_oeb[24]
port 49 nsew signal output
rlabel metal2 s 11794 49200 11850 50000 6 io_oeb[25]
port 50 nsew signal output
rlabel metal2 s 12254 49200 12310 50000 6 io_oeb[26]
port 51 nsew signal output
rlabel metal2 s 12714 49200 12770 50000 6 io_oeb[27]
port 52 nsew signal output
rlabel metal2 s 13174 49200 13230 50000 6 io_oeb[28]
port 53 nsew signal output
rlabel metal2 s 13634 49200 13690 50000 6 io_oeb[29]
port 54 nsew signal output
rlabel metal2 s 1122 49200 1178 50000 6 io_oeb[2]
port 55 nsew signal output
rlabel metal2 s 14094 49200 14150 50000 6 io_oeb[30]
port 56 nsew signal output
rlabel metal2 s 14554 49200 14610 50000 6 io_oeb[31]
port 57 nsew signal output
rlabel metal2 s 1582 49200 1638 50000 6 io_oeb[3]
port 58 nsew signal output
rlabel metal2 s 2042 49200 2098 50000 6 io_oeb[4]
port 59 nsew signal output
rlabel metal2 s 2502 49200 2558 50000 6 io_oeb[5]
port 60 nsew signal output
rlabel metal2 s 2962 49200 3018 50000 6 io_oeb[6]
port 61 nsew signal output
rlabel metal2 s 3422 49200 3478 50000 6 io_oeb[7]
port 62 nsew signal output
rlabel metal2 s 3882 49200 3938 50000 6 io_oeb[8]
port 63 nsew signal output
rlabel metal2 s 4342 49200 4398 50000 6 io_oeb[9]
port 64 nsew signal output
rlabel metal4 s 3910 2128 4230 47376 6 vccd1
port 65 nsew power input
rlabel metal4 s 9840 2128 10160 47376 6 vccd1
port 65 nsew power input
rlabel metal4 s 15771 2128 16091 47376 6 vccd1
port 65 nsew power input
rlabel metal4 s 6874 2128 7194 47376 6 vssd1
port 66 nsew ground input
rlabel metal4 s 12805 2128 13125 47376 6 vssd1
port 66 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 833470
string GDS_FILE /home/salah/AI_CORDIC_LIU/mychip/openlane/cordic/runs/cordic/results/finishing/cordic.magic.gds
string GDS_START 223214
<< end >>


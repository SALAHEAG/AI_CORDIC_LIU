VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cordic
  CLASS BLOCK ;
  FOREIGN cordic ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 246.000 14.630 250.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 246.000 34.870 250.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 246.000 54.650 250.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 28.600 100.000 29.200 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 66.680 100.000 67.280 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 246.000 84.550 250.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 163.240 100.000 163.840 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 221.040 100.000 221.640 ;
    END
  END A[9]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 246.000 4.970 250.000 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 9.560 100.000 10.160 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 246.000 74.430 250.000 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 86.400 100.000 87.000 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 105.440 100.000 106.040 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 182.280 100.000 182.880 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 246.000 94.670 250.000 ;
    END
  END B[9]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END Ci
  PIN Co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END Co
  PIN S[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 246.000 24.750 250.000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 246.000 44.530 250.000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 246.000 64.770 250.000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 47.640 100.000 48.240 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 124.480 100.000 125.080 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 144.200 100.000 144.800 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 202.000 100.000 202.600 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 240.080 100.000 240.680 ;
    END
  END S[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.550 10.640 21.150 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.855 10.640 80.455 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 236.725 ;
      LAYER met1 ;
        RECT 4.670 10.640 94.690 236.880 ;
      LAYER met2 ;
        RECT 5.250 245.720 14.070 246.570 ;
        RECT 14.910 245.720 24.190 246.570 ;
        RECT 25.030 245.720 34.310 246.570 ;
        RECT 35.150 245.720 43.970 246.570 ;
        RECT 44.810 245.720 54.090 246.570 ;
        RECT 54.930 245.720 64.210 246.570 ;
        RECT 65.050 245.720 73.870 246.570 ;
        RECT 74.710 245.720 83.990 246.570 ;
        RECT 84.830 245.720 94.110 246.570 ;
        RECT 4.700 4.280 94.660 245.720 ;
        RECT 4.700 4.000 12.230 4.280 ;
        RECT 13.070 4.000 37.070 4.280 ;
        RECT 37.910 4.000 61.910 4.280 ;
        RECT 62.750 4.000 86.750 4.280 ;
        RECT 87.590 4.000 94.660 4.280 ;
      LAYER met3 ;
        RECT 4.000 239.680 95.600 240.545 ;
        RECT 4.000 225.440 96.000 239.680 ;
        RECT 4.400 224.040 96.000 225.440 ;
        RECT 4.000 222.040 96.000 224.040 ;
        RECT 4.000 220.640 95.600 222.040 ;
        RECT 4.000 203.000 96.000 220.640 ;
        RECT 4.000 201.600 95.600 203.000 ;
        RECT 4.000 183.280 96.000 201.600 ;
        RECT 4.000 181.880 95.600 183.280 ;
        RECT 4.000 175.120 96.000 181.880 ;
        RECT 4.400 173.720 96.000 175.120 ;
        RECT 4.000 164.240 96.000 173.720 ;
        RECT 4.000 162.840 95.600 164.240 ;
        RECT 4.000 145.200 96.000 162.840 ;
        RECT 4.000 143.800 95.600 145.200 ;
        RECT 4.000 125.480 96.000 143.800 ;
        RECT 4.400 124.080 95.600 125.480 ;
        RECT 4.000 106.440 96.000 124.080 ;
        RECT 4.000 105.040 95.600 106.440 ;
        RECT 4.000 87.400 96.000 105.040 ;
        RECT 4.000 86.000 95.600 87.400 ;
        RECT 4.000 75.160 96.000 86.000 ;
        RECT 4.400 73.760 96.000 75.160 ;
        RECT 4.000 67.680 96.000 73.760 ;
        RECT 4.000 66.280 95.600 67.680 ;
        RECT 4.000 48.640 96.000 66.280 ;
        RECT 4.000 47.240 95.600 48.640 ;
        RECT 4.000 29.600 96.000 47.240 ;
        RECT 4.000 28.200 95.600 29.600 ;
        RECT 4.000 25.520 96.000 28.200 ;
        RECT 4.400 24.120 96.000 25.520 ;
        RECT 4.000 10.560 96.000 24.120 ;
        RECT 4.000 9.695 95.600 10.560 ;
      LAYER met4 ;
        RECT 21.550 10.640 33.970 236.880 ;
        RECT 36.370 10.640 48.800 236.880 ;
        RECT 51.200 10.640 63.625 236.880 ;
        RECT 66.025 10.640 78.455 236.880 ;
  END
END cordic
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cordic
  CLASS BLOCK ;
  FOREIGN cordic ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 246.000 73.050 250.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 246.000 81.790 250.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 246.000 85.930 250.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 156.440 100.000 157.040 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 246.000 92.370 250.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 246.000 94.670 250.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 246.000 96.510 250.000 ;
    END
  END A[9]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 31.320 100.000 31.920 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 246.000 77.650 250.000 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 93.880 100.000 94.480 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 246.000 88.230 250.000 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 246.000 98.810 250.000 ;
    END
  END B[9]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 246.000 68.910 250.000 ;
    END
  END Ci
  PIN Co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 246.000 71.210 250.000 ;
    END
  END Co
  PIN S[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 246.000 75.350 250.000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 246.000 79.490 250.000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 246.000 84.090 250.000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 246.000 90.070 250.000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 219.000 100.000 219.600 ;
    END
  END S[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 246.000 1.290 250.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 246.000 22.450 250.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 246.000 24.290 250.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 246.000 26.590 250.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 246.000 28.890 250.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 246.000 30.730 250.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 246.000 33.030 250.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 246.000 34.870 250.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 246.000 37.170 250.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 246.000 39.470 250.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 246.000 41.310 250.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 246.000 3.130 250.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 246.000 43.610 250.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 246.000 45.450 250.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 246.000 47.750 250.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 246.000 50.050 250.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 246.000 51.890 250.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 246.000 54.190 250.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 246.000 56.490 250.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 246.000 58.330 250.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 246.000 60.630 250.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 246.000 62.470 250.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 246.000 5.430 250.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 246.000 64.770 250.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 246.000 67.070 250.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 246.000 7.270 250.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 246.000 9.570 250.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 246.000 11.870 250.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 246.000 13.710 250.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 246.000 16.010 250.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 246.000 17.850 250.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 246.000 20.150 250.000 ;
    END
  END io_oeb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.550 10.640 21.150 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.855 10.640 80.455 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 236.725 ;
      LAYER met1 ;
        RECT 0.070 10.640 98.830 236.880 ;
      LAYER met2 ;
        RECT 0.100 245.720 0.730 246.570 ;
        RECT 1.570 245.720 2.570 246.570 ;
        RECT 3.410 245.720 4.870 246.570 ;
        RECT 5.710 245.720 6.710 246.570 ;
        RECT 7.550 245.720 9.010 246.570 ;
        RECT 9.850 245.720 11.310 246.570 ;
        RECT 12.150 245.720 13.150 246.570 ;
        RECT 13.990 245.720 15.450 246.570 ;
        RECT 16.290 245.720 17.290 246.570 ;
        RECT 18.130 245.720 19.590 246.570 ;
        RECT 20.430 245.720 21.890 246.570 ;
        RECT 22.730 245.720 23.730 246.570 ;
        RECT 24.570 245.720 26.030 246.570 ;
        RECT 26.870 245.720 28.330 246.570 ;
        RECT 29.170 245.720 30.170 246.570 ;
        RECT 31.010 245.720 32.470 246.570 ;
        RECT 33.310 245.720 34.310 246.570 ;
        RECT 35.150 245.720 36.610 246.570 ;
        RECT 37.450 245.720 38.910 246.570 ;
        RECT 39.750 245.720 40.750 246.570 ;
        RECT 41.590 245.720 43.050 246.570 ;
        RECT 43.890 245.720 44.890 246.570 ;
        RECT 45.730 245.720 47.190 246.570 ;
        RECT 48.030 245.720 49.490 246.570 ;
        RECT 50.330 245.720 51.330 246.570 ;
        RECT 52.170 245.720 53.630 246.570 ;
        RECT 54.470 245.720 55.930 246.570 ;
        RECT 56.770 245.720 57.770 246.570 ;
        RECT 58.610 245.720 60.070 246.570 ;
        RECT 60.910 245.720 61.910 246.570 ;
        RECT 62.750 245.720 64.210 246.570 ;
        RECT 65.050 245.720 66.510 246.570 ;
        RECT 67.350 245.720 68.350 246.570 ;
        RECT 69.190 245.720 70.650 246.570 ;
        RECT 71.490 245.720 72.490 246.570 ;
        RECT 73.330 245.720 74.790 246.570 ;
        RECT 75.630 245.720 77.090 246.570 ;
        RECT 77.930 245.720 78.930 246.570 ;
        RECT 79.770 245.720 81.230 246.570 ;
        RECT 82.070 245.720 83.530 246.570 ;
        RECT 84.370 245.720 85.370 246.570 ;
        RECT 86.210 245.720 87.670 246.570 ;
        RECT 88.510 245.720 89.510 246.570 ;
        RECT 90.350 245.720 91.810 246.570 ;
        RECT 92.650 245.720 94.110 246.570 ;
        RECT 94.950 245.720 95.950 246.570 ;
        RECT 96.790 245.720 98.250 246.570 ;
        RECT 0.100 4.280 98.800 245.720 ;
        RECT 0.100 4.000 6.710 4.280 ;
        RECT 7.550 4.000 20.970 4.280 ;
        RECT 21.810 4.000 35.230 4.280 ;
        RECT 36.070 4.000 49.490 4.280 ;
        RECT 50.330 4.000 63.750 4.280 ;
        RECT 64.590 4.000 78.010 4.280 ;
        RECT 78.850 4.000 92.270 4.280 ;
        RECT 93.110 4.000 98.800 4.280 ;
      LAYER met3 ;
        RECT 4.000 229.520 96.000 236.805 ;
        RECT 4.400 228.120 96.000 229.520 ;
        RECT 4.000 220.000 96.000 228.120 ;
        RECT 4.000 218.600 95.600 220.000 ;
        RECT 4.000 188.040 96.000 218.600 ;
        RECT 4.400 186.640 96.000 188.040 ;
        RECT 4.000 157.440 96.000 186.640 ;
        RECT 4.000 156.040 95.600 157.440 ;
        RECT 4.000 146.560 96.000 156.040 ;
        RECT 4.400 145.160 96.000 146.560 ;
        RECT 4.000 104.400 96.000 145.160 ;
        RECT 4.400 103.000 96.000 104.400 ;
        RECT 4.000 94.880 96.000 103.000 ;
        RECT 4.000 93.480 95.600 94.880 ;
        RECT 4.000 62.920 96.000 93.480 ;
        RECT 4.400 61.520 96.000 62.920 ;
        RECT 4.000 32.320 96.000 61.520 ;
        RECT 4.000 30.920 95.600 32.320 ;
        RECT 4.000 21.440 96.000 30.920 ;
        RECT 4.400 20.040 96.000 21.440 ;
        RECT 4.000 10.715 96.000 20.040 ;
      LAYER met4 ;
        RECT 21.550 10.640 33.970 236.880 ;
        RECT 36.370 10.640 48.800 236.880 ;
        RECT 51.200 10.640 63.625 236.880 ;
        RECT 66.025 10.640 78.455 236.880 ;
  END
END cordic
END LIBRARY


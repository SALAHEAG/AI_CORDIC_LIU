VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cordic
  CLASS BLOCK ;
  FOREIGN cordic ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 246.000 82.250 250.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 78.240 100.000 78.840 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 246.000 98.350 250.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 172.080 100.000 172.680 ;
    END
  END A[9]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 246.000 77.650 250.000 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 246.000 79.950 250.000 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 246.000 84.550 250.000 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 109.520 100.000 110.120 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 246.000 91.450 250.000 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 246.000 93.750 250.000 ;
    END
  END B[7]
  PIN B[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 140.800 100.000 141.400 ;
    END
  END B[8]
  PIN B[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 203.360 100.000 203.960 ;
    END
  END B[9]
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 246.000 75.350 250.000 ;
    END
  END Ci
  PIN Co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END Co
  PIN S[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 15.680 100.000 16.280 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 46.960 100.000 47.560 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 246.000 86.850 250.000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 246.000 89.150 250.000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 246.000 96.050 250.000 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 234.640 100.000 235.240 ;
    END
  END S[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 246.000 1.290 250.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 246.000 24.290 250.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 246.000 26.590 250.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 246.000 28.890 250.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 246.000 31.190 250.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 246.000 33.490 250.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 246.000 35.790 250.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 246.000 38.090 250.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 246.000 40.390 250.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 246.000 42.690 250.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 246.000 44.990 250.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 246.000 3.590 250.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 246.000 47.290 250.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 246.000 49.590 250.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 246.000 52.350 250.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 246.000 54.650 250.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 246.000 56.950 250.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 246.000 59.250 250.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 246.000 61.550 250.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 246.000 63.850 250.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 246.000 66.150 250.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 246.000 68.450 250.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 246.000 5.890 250.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 246.000 70.750 250.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 246.000 73.050 250.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 246.000 8.190 250.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 246.000 10.490 250.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 246.000 12.790 250.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 246.000 15.090 250.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 246.000 17.390 250.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 246.000 19.690 250.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 246.000 21.990 250.000 ;
    END
  END io_oeb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.550 10.640 21.150 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.200 10.640 50.800 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.855 10.640 80.455 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 236.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 94.300 236.725 ;
      LAYER met1 ;
        RECT 0.990 10.640 98.370 237.280 ;
      LAYER met2 ;
        RECT 1.570 245.720 3.030 246.570 ;
        RECT 3.870 245.720 5.330 246.570 ;
        RECT 6.170 245.720 7.630 246.570 ;
        RECT 8.470 245.720 9.930 246.570 ;
        RECT 10.770 245.720 12.230 246.570 ;
        RECT 13.070 245.720 14.530 246.570 ;
        RECT 15.370 245.720 16.830 246.570 ;
        RECT 17.670 245.720 19.130 246.570 ;
        RECT 19.970 245.720 21.430 246.570 ;
        RECT 22.270 245.720 23.730 246.570 ;
        RECT 24.570 245.720 26.030 246.570 ;
        RECT 26.870 245.720 28.330 246.570 ;
        RECT 29.170 245.720 30.630 246.570 ;
        RECT 31.470 245.720 32.930 246.570 ;
        RECT 33.770 245.720 35.230 246.570 ;
        RECT 36.070 245.720 37.530 246.570 ;
        RECT 38.370 245.720 39.830 246.570 ;
        RECT 40.670 245.720 42.130 246.570 ;
        RECT 42.970 245.720 44.430 246.570 ;
        RECT 45.270 245.720 46.730 246.570 ;
        RECT 47.570 245.720 49.030 246.570 ;
        RECT 49.870 245.720 51.790 246.570 ;
        RECT 52.630 245.720 54.090 246.570 ;
        RECT 54.930 245.720 56.390 246.570 ;
        RECT 57.230 245.720 58.690 246.570 ;
        RECT 59.530 245.720 60.990 246.570 ;
        RECT 61.830 245.720 63.290 246.570 ;
        RECT 64.130 245.720 65.590 246.570 ;
        RECT 66.430 245.720 67.890 246.570 ;
        RECT 68.730 245.720 70.190 246.570 ;
        RECT 71.030 245.720 72.490 246.570 ;
        RECT 73.330 245.720 74.790 246.570 ;
        RECT 75.630 245.720 77.090 246.570 ;
        RECT 77.930 245.720 79.390 246.570 ;
        RECT 80.230 245.720 81.690 246.570 ;
        RECT 82.530 245.720 83.990 246.570 ;
        RECT 84.830 245.720 86.290 246.570 ;
        RECT 87.130 245.720 88.590 246.570 ;
        RECT 89.430 245.720 90.890 246.570 ;
        RECT 91.730 245.720 93.190 246.570 ;
        RECT 94.030 245.720 95.490 246.570 ;
        RECT 96.330 245.720 97.790 246.570 ;
        RECT 1.020 4.280 98.340 245.720 ;
        RECT 1.020 4.000 12.230 4.280 ;
        RECT 13.070 4.000 37.070 4.280 ;
        RECT 37.910 4.000 61.910 4.280 ;
        RECT 62.750 4.000 86.750 4.280 ;
        RECT 87.590 4.000 98.340 4.280 ;
      LAYER met3 ;
        RECT 4.400 235.640 96.000 236.805 ;
        RECT 4.400 235.600 95.600 235.640 ;
        RECT 4.000 234.240 95.600 235.600 ;
        RECT 4.000 209.120 96.000 234.240 ;
        RECT 4.400 207.720 96.000 209.120 ;
        RECT 4.000 204.360 96.000 207.720 ;
        RECT 4.000 202.960 95.600 204.360 ;
        RECT 4.000 181.240 96.000 202.960 ;
        RECT 4.400 179.840 96.000 181.240 ;
        RECT 4.000 173.080 96.000 179.840 ;
        RECT 4.000 171.680 95.600 173.080 ;
        RECT 4.000 153.360 96.000 171.680 ;
        RECT 4.400 151.960 96.000 153.360 ;
        RECT 4.000 141.800 96.000 151.960 ;
        RECT 4.000 140.400 95.600 141.800 ;
        RECT 4.000 125.480 96.000 140.400 ;
        RECT 4.400 124.080 96.000 125.480 ;
        RECT 4.000 110.520 96.000 124.080 ;
        RECT 4.000 109.120 95.600 110.520 ;
        RECT 4.000 97.600 96.000 109.120 ;
        RECT 4.400 96.200 96.000 97.600 ;
        RECT 4.000 79.240 96.000 96.200 ;
        RECT 4.000 77.840 95.600 79.240 ;
        RECT 4.000 69.720 96.000 77.840 ;
        RECT 4.400 68.320 96.000 69.720 ;
        RECT 4.000 47.960 96.000 68.320 ;
        RECT 4.000 46.560 95.600 47.960 ;
        RECT 4.000 41.840 96.000 46.560 ;
        RECT 4.400 40.440 96.000 41.840 ;
        RECT 4.000 16.680 96.000 40.440 ;
        RECT 4.000 15.280 95.600 16.680 ;
        RECT 4.000 14.640 96.000 15.280 ;
        RECT 4.400 13.240 96.000 14.640 ;
        RECT 4.000 10.715 96.000 13.240 ;
      LAYER met4 ;
        RECT 21.550 10.640 33.970 236.880 ;
        RECT 36.370 10.640 48.800 236.880 ;
        RECT 51.200 10.640 63.625 236.880 ;
        RECT 66.025 10.640 78.455 236.880 ;
        RECT 80.855 10.640 83.425 236.880 ;
  END
END cordic
END LIBRARY

